`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/10/2019 07:18:43 PM
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(
input wire clk,
input wire reset,
input wire clk_enable,
input wire [7:0] pixelL_in,
input wire [7:0] pixelR_in,
output ce_out,
output en2,
output [7:0] pixel_out
);

wire [7:0] rowL_0;
wire [7:0] rowL_1;
wire [7:0] rowL_2;
wire [7:0] rowL_3;
wire [7:0] rowL_4;
wire [7:0] rowL_5;
wire [7:0] rowL_6;
wire [7:0] rowL_7;
wire [7:0] rowL_8;
wire [7:0] rowL_9;
wire [7:0] rowL_10;
wire [7:0] rowL_11;
wire [7:0] rowL_12;
wire [7:0] rowL_13;
wire [7:0] rowL_14;
wire [7:0] rowL_15;
wire [7:0] rowL_16;
wire [7:0] rowL_17;
wire [7:0] rowL_18;
wire [7:0] rowL_19;
wire [7:0] rowL_20;
wire [7:0] rowL_21;
wire [7:0] rowL_22;
wire [7:0] rowL_23;
wire [7:0] rowL_24;
wire [7:0] rowL_25;
wire [7:0] rowL_26;
wire [7:0] rowL_27;
wire [7:0] rowL_28;
wire [7:0] rowL_29;
wire [7:0] rowL_30;
wire [7:0] rowL_31;
wire [7:0] rowL_32;
wire [7:0] rowL_33;
wire [7:0] rowL_34;
wire [7:0] rowL_35;
wire [7:0] rowL_36;
wire [7:0] rowL_37;
wire [7:0] rowL_38;
wire [7:0] rowL_39;
wire [7:0] rowL_40;
wire [7:0] rowL_41;
wire [7:0] rowL_42;
wire [7:0] rowL_43;
wire [7:0] rowL_44;
wire [7:0] rowL_45;
wire [7:0] rowL_46;
wire [7:0] rowL_47;
wire [7:0] rowL_48;
wire [7:0] rowL_49;
wire [7:0] rowL_50;
wire [7:0] rowL_51;
wire [7:0] rowL_52;
wire [7:0] rowL_53;
wire [7:0] rowL_54;
wire [7:0] rowL_55;
wire [7:0] rowL_56;
wire [7:0] rowL_57;
wire [7:0] rowL_58;
wire [7:0] rowL_59;
wire [7:0] rowL_60;
wire [7:0] rowL_61;
wire [7:0] rowL_62;
wire [7:0] rowL_63;
wire [7:0] rowL_64;
wire [7:0] rowL_65;
wire [7:0] rowL_66;
wire [7:0] rowL_67;
wire [7:0] rowL_68;
wire [7:0] rowL_69;
wire [7:0] rowL_70;
wire [7:0] rowL_71;
wire [7:0] rowL_72;
wire [7:0] rowL_73;
wire [7:0] rowL_74;
wire [7:0] rowL_75;
wire [7:0] rowL_76;
wire [7:0] rowL_77;
wire [7:0] rowL_78;
wire [7:0] rowL_79;
wire [7:0] rowL_80;
wire [7:0] rowL_81;
wire [7:0] rowL_82;
wire [7:0] rowL_83;
wire [7:0] rowL_84;
wire [7:0] rowL_85;
wire [7:0] rowL_86;
wire [7:0] rowL_87;
wire [7:0] rowL_88;
wire [7:0] rowL_89;
wire [7:0] rowL_90;
wire [7:0] rowL_91;
wire [7:0] rowL_92;
wire [7:0] rowL_93;
wire [7:0] rowL_94;
wire [7:0] rowL_95;
wire [7:0] rowL_96;
wire [7:0] rowL_97;
wire [7:0] rowL_98;
wire [7:0] rowL_99;
wire [7:0] rowL_100;
wire [7:0] rowL_101;
wire [7:0] rowL_102;
wire [7:0] rowL_103;
wire [7:0] rowL_104;
wire [7:0] rowL_105;
wire [7:0] rowL_106;
wire [7:0] rowL_107;
wire [7:0] rowL_108;
wire [7:0] rowL_109;
wire [7:0] rowL_110;
wire [7:0] rowL_111;
wire [7:0] rowL_112;
wire [7:0] rowL_113;
wire [7:0] rowL_114;
wire [7:0] rowL_115;
wire [7:0] rowL_116;
wire [7:0] rowL_117;
wire [7:0] rowL_118;
wire [7:0] rowL_119;
wire [7:0] rowL_120;
wire [7:0] rowL_121;
wire [7:0] rowL_122;
wire [7:0] rowL_123;
wire [7:0] rowL_124;
wire [7:0] rowL_125;
wire [7:0] rowL_126;
wire [7:0] rowL_127;
wire [7:0] rowL_128;
wire [7:0] rowL_129;
wire [7:0] rowL_130;
wire [7:0] rowL_131;
wire [7:0] rowL_132;
wire [7:0] rowL_133;
wire [7:0] rowL_134;
wire [7:0] rowL_135;
wire [7:0] rowL_136;
wire [7:0] rowL_137;
wire [7:0] rowL_138;
wire [7:0] rowL_139;
wire [7:0] rowL_140;
wire [7:0] rowL_141;
wire [7:0] rowL_142;
wire [7:0] rowL_143;
wire [7:0] rowL_144;
wire [7:0] rowL_145;
wire [7:0] rowL_146;
wire [7:0] rowL_147;
wire [7:0] rowL_148;
wire [7:0] rowL_149;
wire [7:0] rowL_150;
wire [7:0] rowL_151;
wire [7:0] rowL_152;
wire [7:0] rowL_153;
wire [7:0] rowL_154;
wire [7:0] rowL_155;
wire [7:0] rowL_156;
wire [7:0] rowL_157;
wire [7:0] rowL_158;
wire [7:0] rowL_159;
wire [7:0] rowL_160;
wire [7:0] rowL_161;
wire [7:0] rowL_162;
wire [7:0] rowL_163;
wire [7:0] rowL_164;
wire [7:0] rowL_165;
wire [7:0] rowL_166;
wire [7:0] rowL_167;
wire [7:0] rowL_168;
wire [7:0] rowL_169;
wire [7:0] rowL_170;
wire [7:0] rowL_171;
wire [7:0] rowL_172;
wire [7:0] rowL_173;
wire [7:0] rowL_174;
wire [7:0] rowL_175;
wire [7:0] rowL_176;
wire [7:0] rowL_177;
wire [7:0] rowL_178;
wire [7:0] rowL_179;
wire [7:0] rowL_180;
wire [7:0] rowL_181;
wire [7:0] rowL_182;
wire [7:0] rowL_183;
wire [7:0] rowL_184;
wire [7:0] rowL_185;
wire [7:0] rowL_186;
wire [7:0] rowL_187;
wire [7:0] rowL_188;
wire [7:0] rowL_189;
wire [7:0] rowL_190;
wire [7:0] rowL_191;
wire [7:0] rowL_192;
wire [7:0] rowL_193;
wire [7:0] rowL_194;
wire [7:0] rowL_195;
wire [7:0] rowL_196;
wire [7:0] rowL_197;
wire [7:0] rowL_198;
wire [7:0] rowL_199;
wire [7:0] rowL_200;
wire [7:0] rowL_201;
wire [7:0] rowL_202;
wire [7:0] rowL_203;
wire [7:0] rowL_204;
wire [7:0] rowL_205;
wire [7:0] rowL_206;
wire [7:0] rowL_207;
wire [7:0] rowL_208;
wire [7:0] rowL_209;
wire [7:0] rowL_210;
wire [7:0] rowL_211;
wire [7:0] rowL_212;
wire [7:0] rowL_213;
wire [7:0] rowL_214;
wire [7:0] rowL_215;
wire [7:0] rowL_216;
wire [7:0] rowL_217;
wire [7:0] rowL_218;
wire [7:0] rowL_219;
wire [7:0] rowL_220;
wire [7:0] rowL_221;
wire [7:0] rowL_222;
wire [7:0] rowL_223;
wire [7:0] rowL_224;
wire [7:0] rowL_225;
wire [7:0] rowL_226;
wire [7:0] rowL_227;
wire [7:0] rowL_228;
wire [7:0] rowL_229;
wire [7:0] rowL_230;
wire [7:0] rowL_231;
wire [7:0] rowL_232;
wire [7:0] rowL_233;
wire [7:0] rowL_234;
wire [7:0] rowL_235;
wire [7:0] rowL_236;
wire [7:0] rowL_237;
wire [7:0] rowL_238;
wire [7:0] rowL_239;
wire [7:0] rowL_240;
wire [7:0] rowL_241;
wire [7:0] rowL_242;
wire [7:0] rowL_243;
wire [7:0] rowL_244;
wire [7:0] rowL_245;
wire [7:0] rowL_246;
wire [7:0] rowL_247;
wire [7:0] rowL_248;
wire [7:0] rowL_249;
wire [7:0] rowL_250;
wire [7:0] rowL_251;
wire [7:0] rowL_252;
wire [7:0] rowL_253;
wire [7:0] rowL_254;
wire [7:0] rowL_255;
wire [7:0] rowL_256;
wire [7:0] rowL_257;
wire [7:0] rowL_258;
wire [7:0] rowL_259;
wire [7:0] rowL_260;
wire [7:0] rowL_261;
wire [7:0] rowL_262;
wire [7:0] rowL_263;
wire [7:0] rowL_264;
wire [7:0] rowL_265;
wire [7:0] rowL_266;
wire [7:0] rowL_267;
wire [7:0] rowL_268;
wire [7:0] rowL_269;
wire [7:0] rowL_270;
wire [7:0] rowL_271;
wire [7:0] rowL_272;
wire [7:0] rowL_273;
wire [7:0] rowL_274;
wire [7:0] rowL_275;
wire [7:0] rowL_276;
wire [7:0] rowL_277;
wire [7:0] rowL_278;
wire [7:0] rowL_279;
wire [7:0] rowL_280;
wire [7:0] rowL_281;
wire [7:0] rowL_282;
wire [7:0] rowL_283;
wire [7:0] rowL_284;
wire [7:0] rowL_285;
wire [7:0] rowL_286;
wire [7:0] rowL_287;
wire [7:0] rowL_288;
wire [7:0] rowL_289;
wire [7:0] rowL_290;
wire [7:0] rowL_291;
wire [7:0] rowL_292;
wire [7:0] rowL_293;
wire [7:0] rowL_294;
wire [7:0] rowL_295;
wire [7:0] rowL_296;
wire [7:0] rowL_297;
wire [7:0] rowL_298;
wire [7:0] rowL_299;
wire [7:0] rowL_300;
wire [7:0] rowL_301;
wire [7:0] rowL_302;
wire [7:0] rowL_303;
wire [7:0] rowL_304;
wire [7:0] rowL_305;
wire [7:0] rowL_306;
wire [7:0] rowL_307;
wire [7:0] rowL_308;
wire [7:0] rowL_309;
wire [7:0] rowL_310;
wire [7:0] rowL_311;
wire [7:0] rowL_312;
wire [7:0] rowL_313;
wire [7:0] rowL_314;
wire [7:0] rowL_315;
wire [7:0] rowL_316;
wire [7:0] rowL_317;
wire [7:0] rowL_318;
wire [7:0] rowL_319;
wire [7:0] rowL_320;
wire [7:0] rowL_321;
wire [7:0] rowL_322;
wire [7:0] rowL_323;
wire [7:0] rowL_324;
wire [7:0] rowL_325;
wire [7:0] rowL_326;
wire [7:0] rowL_327;
wire [7:0] rowL_328;
wire [7:0] rowL_329;
wire [7:0] rowL_330;
wire [7:0] rowL_331;
wire [7:0] rowL_332;
wire [7:0] rowL_333;
wire [7:0] rowL_334;
wire [7:0] rowL_335;
wire [7:0] rowL_336;
wire [7:0] rowL_337;
wire [7:0] rowL_338;
wire [7:0] rowL_339;
wire [7:0] rowL_340;
wire [7:0] rowL_341;
wire [7:0] rowL_342;
wire [7:0] rowL_343;
wire [7:0] rowL_344;
wire [7:0] rowL_345;
wire [7:0] rowL_346;
wire [7:0] rowL_347;
wire [7:0] rowL_348;
wire [7:0] rowL_349;
wire [7:0] rowL_350;
wire [7:0] rowL_351;
wire [7:0] rowL_352;
wire [7:0] rowL_353;
wire [7:0] rowL_354;
wire [7:0] rowL_355;
wire [7:0] rowL_356;
wire [7:0] rowL_357;
wire [7:0] rowL_358;
wire [7:0] rowL_359;
wire [7:0] rowL_360;
wire [7:0] rowL_361;
wire [7:0] rowL_362;
wire [7:0] rowL_363;
wire [7:0] rowL_364;
wire [7:0] rowL_365;
wire [7:0] rowL_366;
wire [7:0] rowL_367;
wire [7:0] rowL_368;
wire [7:0] rowL_369;
wire [7:0] rowL_370;
wire [7:0] rowL_371;
wire [7:0] rowL_372;
wire [7:0] rowL_373;
wire [7:0] rowL_374;
wire [7:0] rowL_375;
wire [7:0] rowL_376;
wire [7:0] rowL_377;
wire [7:0] rowL_378;
wire [7:0] rowL_379;
wire [7:0] rowL_380;
wire [7:0] rowL_381;
wire [7:0] rowL_382;
wire [7:0] rowL_383;
wire [7:0] rowL_384;
wire [7:0] rowL_385;
wire [7:0] rowL_386;
wire [7:0] rowL_387;
wire [7:0] rowL_388;
wire [7:0] rowL_389;
wire [7:0] rowL_390;
wire [7:0] rowL_391;
wire [7:0] rowL_392;
wire [7:0] rowL_393;
wire [7:0] rowL_394;
wire [7:0] rowL_395;
wire [7:0] rowL_396;
wire [7:0] rowL_397;
wire [7:0] rowL_398;
wire [7:0] rowL_399;
wire [7:0] rowL_400;
wire [7:0] rowL_401;
wire [7:0] rowL_402;
wire [7:0] rowL_403;
wire [7:0] rowL_404;
wire [7:0] rowL_405;
wire [7:0] rowL_406;
wire [7:0] rowL_407;
wire [7:0] rowL_408;
wire [7:0] rowL_409;
wire [7:0] rowL_410;
wire [7:0] rowL_411;
wire [7:0] rowL_412;
wire [7:0] rowL_413;
wire [7:0] rowL_414;
wire [7:0] rowL_415;
wire [7:0] rowL_416;
wire [7:0] rowL_417;
wire [7:0] rowL_418;
wire [7:0] rowL_419;
wire [7:0] rowL_420;
wire [7:0] rowL_421;
wire [7:0] rowL_422;
wire [7:0] rowL_423;
wire [7:0] rowL_424;
wire [7:0] rowL_425;
wire [7:0] rowL_426;
wire [7:0] rowL_427;
wire [7:0] rowL_428;
wire [7:0] rowL_429;
wire [7:0] rowL_430;
wire [7:0] rowL_431;
wire [7:0] rowL_432;
wire [7:0] rowL_433;
wire [7:0] rowL_434;
wire [7:0] rowL_435;
wire [7:0] rowL_436;
wire [7:0] rowL_437;
wire [7:0] rowL_438;
wire [7:0] rowL_439;
wire [7:0] rowL_440;
wire [7:0] rowL_441;
wire [7:0] rowL_442;
wire [7:0] rowL_443;
wire [7:0] rowL_444;
wire [7:0] rowL_445;
wire [7:0] rowL_446;
wire [7:0] rowL_447;
wire [7:0] rowL_448;
wire [7:0] rowL_449;
wire [7:0] rowL_450;
wire [7:0] rowL_451;
wire [7:0] rowL_452;
wire [7:0] rowL_453;
wire [7:0] rowL_454;
wire [7:0] rowL_455;
wire [7:0] rowL_456;
wire [7:0] rowL_457;
wire [7:0] rowL_458;
wire [7:0] rowL_459;
wire [7:0] rowL_460;
wire [7:0] rowL_461;
wire [7:0] rowL_462;
wire [7:0] rowL_463;
wire [7:0] rowL_464;
wire [7:0] rowL_465;
wire [7:0] rowL_466;
wire [7:0] rowL_467;
wire [7:0] rowL_468;
wire [7:0] rowL_469;
wire [7:0] rowL_470;
wire [7:0] rowL_471;
wire [7:0] rowL_472;
wire [7:0] rowL_473;
wire [7:0] rowL_474;
wire [7:0] rowL_475;
wire [7:0] rowL_476;
wire [7:0] rowL_477;
wire [7:0] rowL_478;
wire [7:0] rowL_479;
wire [7:0] rowL_480;
wire [7:0] rowL_481;
wire [7:0] rowL_482;
wire [7:0] rowL_483;
wire [7:0] rowL_484;
wire [7:0] rowL_485;
wire [7:0] rowL_486;
wire [7:0] rowL_487;
wire [7:0] rowL_488;
wire [7:0] rowL_489;
wire [7:0] rowL_490;
wire [7:0] rowL_491;
wire [7:0] rowL_492;
wire [7:0] rowL_493;
wire [7:0] rowL_494;
wire [7:0] rowL_495;
wire [7:0] rowL_496;
wire [7:0] rowL_497;
wire [7:0] rowL_498;
wire [7:0] rowL_499;
wire [7:0] rowL_500;
wire [7:0] rowL_501;
wire [7:0] rowL_502;
wire [7:0] rowL_503;
wire [7:0] rowL_504;
wire [7:0] rowL_505;
wire [7:0] rowL_506;
wire [7:0] rowL_507;
wire [7:0] rowL_508;
wire [7:0] rowL_509;
wire [7:0] rowL_510;
wire [7:0] rowL_511;
wire [7:0] rowL_512;
wire [7:0] rowL_513;
wire [7:0] rowL_514;
wire [7:0] rowL_515;
wire [7:0] rowL_516;
wire [7:0] rowL_517;
wire [7:0] rowL_518;
wire [7:0] rowL_519;
wire [7:0] rowL_520;
wire [7:0] rowL_521;
wire [7:0] rowL_522;
wire [7:0] rowL_523;
wire [7:0] rowL_524;
wire [7:0] rowL_525;
wire [7:0] rowL_526;
wire [7:0] rowL_527;
wire [7:0] rowL_528;
wire [7:0] rowL_529;
wire [7:0] rowL_530;
wire [7:0] rowL_531;
wire [7:0] rowL_532;
wire [7:0] rowL_533;
wire [7:0] rowL_534;
wire [7:0] rowL_535;
wire [7:0] rowL_536;
wire [7:0] rowL_537;
wire [7:0] rowL_538;
wire [7:0] rowL_539;
wire [7:0] rowL_540;
wire [7:0] rowL_541;
wire [7:0] rowL_542;
wire [7:0] rowL_543;
wire [7:0] rowL_544;
wire [7:0] rowL_545;
wire [7:0] rowL_546;
wire [7:0] rowL_547;
wire [7:0] rowL_548;
wire [7:0] rowL_549;
wire [7:0] rowL_550;
wire [7:0] rowL_551;
wire [7:0] rowL_552;
wire [7:0] rowL_553;
wire [7:0] rowL_554;
wire [7:0] rowL_555;
wire [7:0] rowL_556;
wire [7:0] rowL_557;
wire [7:0] rowL_558;
wire [7:0] rowL_559;
wire [7:0] rowL_560;
wire [7:0] rowL_561;
wire [7:0] rowL_562;
wire [7:0] rowL_563;
wire [7:0] rowL_564;
wire [7:0] rowL_565;
wire [7:0] rowL_566;
wire [7:0] rowL_567;
wire [7:0] rowL_568;
wire [7:0] rowL_569;
wire [7:0] rowL_570;
wire [7:0] rowL_571;
wire [7:0] rowL_572;
wire [7:0] rowL_573;
wire [7:0] rowL_574;
wire [7:0] rowL_575;
wire [7:0] rowL_576;
wire [7:0] rowL_577;
wire [7:0] rowL_578;
wire [7:0] rowL_579;
wire [7:0] rowL_580;
wire [7:0] rowL_581;
wire [7:0] rowL_582;
wire [7:0] rowL_583;
wire [7:0] rowL_584;
wire [7:0] rowL_585;
wire [7:0] rowL_586;
wire [7:0] rowL_587;
wire [7:0] rowL_588;
wire [7:0] rowL_589;
wire [7:0] rowL_590;
wire [7:0] rowL_591;
wire [7:0] rowL_592;
wire [7:0] rowL_593;
wire [7:0] rowL_594;
wire [7:0] rowL_595;
wire [7:0] rowL_596;
wire [7:0] rowL_597;
wire [7:0] rowL_598;
wire [7:0] rowL_599;
wire [7:0] rowL_600;
wire [7:0] rowL_601;
wire [7:0] rowL_602;
wire [7:0] rowL_603;
wire [7:0] rowL_604;
wire [7:0] rowL_605;
wire [7:0] rowL_606;
wire [7:0] rowL_607;
wire [7:0] rowL_608;
wire [7:0] rowL_609;
wire [7:0] rowL_610;
wire [7:0] rowL_611;
wire [7:0] rowL_612;
wire [7:0] rowL_613;
wire [7:0] rowL_614;
wire [7:0] rowL_615;
wire [7:0] rowL_616;
wire [7:0] rowL_617;
wire [7:0] rowL_618;
wire [7:0] rowL_619;
wire [7:0] rowL_620;
wire [7:0] rowL_621;
wire [7:0] rowL_622;
wire [7:0] rowL_623;
wire [7:0] rowL_624;
wire [7:0] rowL_625;
wire [7:0] rowL_626;
wire [7:0] rowL_627;
wire [7:0] rowL_628;
wire [7:0] rowL_629;
wire [7:0] rowL_630;
wire [7:0] rowL_631;
wire [7:0] rowL_632;
wire [7:0] rowL_633;
wire [7:0] rowL_634;
wire [7:0] rowL_635;
wire [7:0] rowL_636;
wire [7:0] rowL_637;
wire [7:0] rowL_638;
wire [7:0] rowL_639;

wire [7:0] rowR_0;
wire [7:0] rowR_1;
wire [7:0] rowR_2;
wire [7:0] rowR_3;
wire [7:0] rowR_4;
wire [7:0] rowR_5;
wire [7:0] rowR_6;
wire [7:0] rowR_7;
wire [7:0] rowR_8;
wire [7:0] rowR_9;
wire [7:0] rowR_10;
wire [7:0] rowR_11;
wire [7:0] rowR_12;
wire [7:0] rowR_13;
wire [7:0] rowR_14;
wire [7:0] rowR_15;
wire [7:0] rowR_16;
wire [7:0] rowR_17;
wire [7:0] rowR_18;
wire [7:0] rowR_19;
wire [7:0] rowR_20;
wire [7:0] rowR_21;
wire [7:0] rowR_22;
wire [7:0] rowR_23;
wire [7:0] rowR_24;
wire [7:0] rowR_25;
wire [7:0] rowR_26;
wire [7:0] rowR_27;
wire [7:0] rowR_28;
wire [7:0] rowR_29;
wire [7:0] rowR_30;
wire [7:0] rowR_31;
wire [7:0] rowR_32;
wire [7:0] rowR_33;
wire [7:0] rowR_34;
wire [7:0] rowR_35;
wire [7:0] rowR_36;
wire [7:0] rowR_37;
wire [7:0] rowR_38;
wire [7:0] rowR_39;
wire [7:0] rowR_40;
wire [7:0] rowR_41;
wire [7:0] rowR_42;
wire [7:0] rowR_43;
wire [7:0] rowR_44;
wire [7:0] rowR_45;
wire [7:0] rowR_46;
wire [7:0] rowR_47;
wire [7:0] rowR_48;
wire [7:0] rowR_49;
wire [7:0] rowR_50;
wire [7:0] rowR_51;
wire [7:0] rowR_52;
wire [7:0] rowR_53;
wire [7:0] rowR_54;
wire [7:0] rowR_55;
wire [7:0] rowR_56;
wire [7:0] rowR_57;
wire [7:0] rowR_58;
wire [7:0] rowR_59;
wire [7:0] rowR_60;
wire [7:0] rowR_61;
wire [7:0] rowR_62;
wire [7:0] rowR_63;
wire [7:0] rowR_64;
wire [7:0] rowR_65;
wire [7:0] rowR_66;
wire [7:0] rowR_67;
wire [7:0] rowR_68;
wire [7:0] rowR_69;
wire [7:0] rowR_70;
wire [7:0] rowR_71;
wire [7:0] rowR_72;
wire [7:0] rowR_73;
wire [7:0] rowR_74;
wire [7:0] rowR_75;
wire [7:0] rowR_76;
wire [7:0] rowR_77;
wire [7:0] rowR_78;
wire [7:0] rowR_79;
wire [7:0] rowR_80;
wire [7:0] rowR_81;
wire [7:0] rowR_82;
wire [7:0] rowR_83;
wire [7:0] rowR_84;
wire [7:0] rowR_85;
wire [7:0] rowR_86;
wire [7:0] rowR_87;
wire [7:0] rowR_88;
wire [7:0] rowR_89;
wire [7:0] rowR_90;
wire [7:0] rowR_91;
wire [7:0] rowR_92;
wire [7:0] rowR_93;
wire [7:0] rowR_94;
wire [7:0] rowR_95;
wire [7:0] rowR_96;
wire [7:0] rowR_97;
wire [7:0] rowR_98;
wire [7:0] rowR_99;
wire [7:0] rowR_100;
wire [7:0] rowR_101;
wire [7:0] rowR_102;
wire [7:0] rowR_103;
wire [7:0] rowR_104;
wire [7:0] rowR_105;
wire [7:0] rowR_106;
wire [7:0] rowR_107;
wire [7:0] rowR_108;
wire [7:0] rowR_109;
wire [7:0] rowR_110;
wire [7:0] rowR_111;
wire [7:0] rowR_112;
wire [7:0] rowR_113;
wire [7:0] rowR_114;
wire [7:0] rowR_115;
wire [7:0] rowR_116;
wire [7:0] rowR_117;
wire [7:0] rowR_118;
wire [7:0] rowR_119;
wire [7:0] rowR_120;
wire [7:0] rowR_121;
wire [7:0] rowR_122;
wire [7:0] rowR_123;
wire [7:0] rowR_124;
wire [7:0] rowR_125;
wire [7:0] rowR_126;
wire [7:0] rowR_127;
wire [7:0] rowR_128;
wire [7:0] rowR_129;
wire [7:0] rowR_130;
wire [7:0] rowR_131;
wire [7:0] rowR_132;
wire [7:0] rowR_133;
wire [7:0] rowR_134;
wire [7:0] rowR_135;
wire [7:0] rowR_136;
wire [7:0] rowR_137;
wire [7:0] rowR_138;
wire [7:0] rowR_139;
wire [7:0] rowR_140;
wire [7:0] rowR_141;
wire [7:0] rowR_142;
wire [7:0] rowR_143;
wire [7:0] rowR_144;
wire [7:0] rowR_145;
wire [7:0] rowR_146;
wire [7:0] rowR_147;
wire [7:0] rowR_148;
wire [7:0] rowR_149;
wire [7:0] rowR_150;
wire [7:0] rowR_151;
wire [7:0] rowR_152;
wire [7:0] rowR_153;
wire [7:0] rowR_154;
wire [7:0] rowR_155;
wire [7:0] rowR_156;
wire [7:0] rowR_157;
wire [7:0] rowR_158;
wire [7:0] rowR_159;
wire [7:0] rowR_160;
wire [7:0] rowR_161;
wire [7:0] rowR_162;
wire [7:0] rowR_163;
wire [7:0] rowR_164;
wire [7:0] rowR_165;
wire [7:0] rowR_166;
wire [7:0] rowR_167;
wire [7:0] rowR_168;
wire [7:0] rowR_169;
wire [7:0] rowR_170;
wire [7:0] rowR_171;
wire [7:0] rowR_172;
wire [7:0] rowR_173;
wire [7:0] rowR_174;
wire [7:0] rowR_175;
wire [7:0] rowR_176;
wire [7:0] rowR_177;
wire [7:0] rowR_178;
wire [7:0] rowR_179;
wire [7:0] rowR_180;
wire [7:0] rowR_181;
wire [7:0] rowR_182;
wire [7:0] rowR_183;
wire [7:0] rowR_184;
wire [7:0] rowR_185;
wire [7:0] rowR_186;
wire [7:0] rowR_187;
wire [7:0] rowR_188;
wire [7:0] rowR_189;
wire [7:0] rowR_190;
wire [7:0] rowR_191;
wire [7:0] rowR_192;
wire [7:0] rowR_193;
wire [7:0] rowR_194;
wire [7:0] rowR_195;
wire [7:0] rowR_196;
wire [7:0] rowR_197;
wire [7:0] rowR_198;
wire [7:0] rowR_199;
wire [7:0] rowR_200;
wire [7:0] rowR_201;
wire [7:0] rowR_202;
wire [7:0] rowR_203;
wire [7:0] rowR_204;
wire [7:0] rowR_205;
wire [7:0] rowR_206;
wire [7:0] rowR_207;
wire [7:0] rowR_208;
wire [7:0] rowR_209;
wire [7:0] rowR_210;
wire [7:0] rowR_211;
wire [7:0] rowR_212;
wire [7:0] rowR_213;
wire [7:0] rowR_214;
wire [7:0] rowR_215;
wire [7:0] rowR_216;
wire [7:0] rowR_217;
wire [7:0] rowR_218;
wire [7:0] rowR_219;
wire [7:0] rowR_220;
wire [7:0] rowR_221;
wire [7:0] rowR_222;
wire [7:0] rowR_223;
wire [7:0] rowR_224;
wire [7:0] rowR_225;
wire [7:0] rowR_226;
wire [7:0] rowR_227;
wire [7:0] rowR_228;
wire [7:0] rowR_229;
wire [7:0] rowR_230;
wire [7:0] rowR_231;
wire [7:0] rowR_232;
wire [7:0] rowR_233;
wire [7:0] rowR_234;
wire [7:0] rowR_235;
wire [7:0] rowR_236;
wire [7:0] rowR_237;
wire [7:0] rowR_238;
wire [7:0] rowR_239;
wire [7:0] rowR_240;
wire [7:0] rowR_241;
wire [7:0] rowR_242;
wire [7:0] rowR_243;
wire [7:0] rowR_244;
wire [7:0] rowR_245;
wire [7:0] rowR_246;
wire [7:0] rowR_247;
wire [7:0] rowR_248;
wire [7:0] rowR_249;
wire [7:0] rowR_250;
wire [7:0] rowR_251;
wire [7:0] rowR_252;
wire [7:0] rowR_253;
wire [7:0] rowR_254;
wire [7:0] rowR_255;
wire [7:0] rowR_256;
wire [7:0] rowR_257;
wire [7:0] rowR_258;
wire [7:0] rowR_259;
wire [7:0] rowR_260;
wire [7:0] rowR_261;
wire [7:0] rowR_262;
wire [7:0] rowR_263;
wire [7:0] rowR_264;
wire [7:0] rowR_265;
wire [7:0] rowR_266;
wire [7:0] rowR_267;
wire [7:0] rowR_268;
wire [7:0] rowR_269;
wire [7:0] rowR_270;
wire [7:0] rowR_271;
wire [7:0] rowR_272;
wire [7:0] rowR_273;
wire [7:0] rowR_274;
wire [7:0] rowR_275;
wire [7:0] rowR_276;
wire [7:0] rowR_277;
wire [7:0] rowR_278;
wire [7:0] rowR_279;
wire [7:0] rowR_280;
wire [7:0] rowR_281;
wire [7:0] rowR_282;
wire [7:0] rowR_283;
wire [7:0] rowR_284;
wire [7:0] rowR_285;
wire [7:0] rowR_286;
wire [7:0] rowR_287;
wire [7:0] rowR_288;
wire [7:0] rowR_289;
wire [7:0] rowR_290;
wire [7:0] rowR_291;
wire [7:0] rowR_292;
wire [7:0] rowR_293;
wire [7:0] rowR_294;
wire [7:0] rowR_295;
wire [7:0] rowR_296;
wire [7:0] rowR_297;
wire [7:0] rowR_298;
wire [7:0] rowR_299;
wire [7:0] rowR_300;
wire [7:0] rowR_301;
wire [7:0] rowR_302;
wire [7:0] rowR_303;
wire [7:0] rowR_304;
wire [7:0] rowR_305;
wire [7:0] rowR_306;
wire [7:0] rowR_307;
wire [7:0] rowR_308;
wire [7:0] rowR_309;
wire [7:0] rowR_310;
wire [7:0] rowR_311;
wire [7:0] rowR_312;
wire [7:0] rowR_313;
wire [7:0] rowR_314;
wire [7:0] rowR_315;
wire [7:0] rowR_316;
wire [7:0] rowR_317;
wire [7:0] rowR_318;
wire [7:0] rowR_319;
wire [7:0] rowR_320;
wire [7:0] rowR_321;
wire [7:0] rowR_322;
wire [7:0] rowR_323;
wire [7:0] rowR_324;
wire [7:0] rowR_325;
wire [7:0] rowR_326;
wire [7:0] rowR_327;
wire [7:0] rowR_328;
wire [7:0] rowR_329;
wire [7:0] rowR_330;
wire [7:0] rowR_331;
wire [7:0] rowR_332;
wire [7:0] rowR_333;
wire [7:0] rowR_334;
wire [7:0] rowR_335;
wire [7:0] rowR_336;
wire [7:0] rowR_337;
wire [7:0] rowR_338;
wire [7:0] rowR_339;
wire [7:0] rowR_340;
wire [7:0] rowR_341;
wire [7:0] rowR_342;
wire [7:0] rowR_343;
wire [7:0] rowR_344;
wire [7:0] rowR_345;
wire [7:0] rowR_346;
wire [7:0] rowR_347;
wire [7:0] rowR_348;
wire [7:0] rowR_349;
wire [7:0] rowR_350;
wire [7:0] rowR_351;
wire [7:0] rowR_352;
wire [7:0] rowR_353;
wire [7:0] rowR_354;
wire [7:0] rowR_355;
wire [7:0] rowR_356;
wire [7:0] rowR_357;
wire [7:0] rowR_358;
wire [7:0] rowR_359;
wire [7:0] rowR_360;
wire [7:0] rowR_361;
wire [7:0] rowR_362;
wire [7:0] rowR_363;
wire [7:0] rowR_364;
wire [7:0] rowR_365;
wire [7:0] rowR_366;
wire [7:0] rowR_367;
wire [7:0] rowR_368;
wire [7:0] rowR_369;
wire [7:0] rowR_370;
wire [7:0] rowR_371;
wire [7:0] rowR_372;
wire [7:0] rowR_373;
wire [7:0] rowR_374;
wire [7:0] rowR_375;
wire [7:0] rowR_376;
wire [7:0] rowR_377;
wire [7:0] rowR_378;
wire [7:0] rowR_379;
wire [7:0] rowR_380;
wire [7:0] rowR_381;
wire [7:0] rowR_382;
wire [7:0] rowR_383;
wire [7:0] rowR_384;
wire [7:0] rowR_385;
wire [7:0] rowR_386;
wire [7:0] rowR_387;
wire [7:0] rowR_388;
wire [7:0] rowR_389;
wire [7:0] rowR_390;
wire [7:0] rowR_391;
wire [7:0] rowR_392;
wire [7:0] rowR_393;
wire [7:0] rowR_394;
wire [7:0] rowR_395;
wire [7:0] rowR_396;
wire [7:0] rowR_397;
wire [7:0] rowR_398;
wire [7:0] rowR_399;
wire [7:0] rowR_400;
wire [7:0] rowR_401;
wire [7:0] rowR_402;
wire [7:0] rowR_403;
wire [7:0] rowR_404;
wire [7:0] rowR_405;
wire [7:0] rowR_406;
wire [7:0] rowR_407;
wire [7:0] rowR_408;
wire [7:0] rowR_409;
wire [7:0] rowR_410;
wire [7:0] rowR_411;
wire [7:0] rowR_412;
wire [7:0] rowR_413;
wire [7:0] rowR_414;
wire [7:0] rowR_415;
wire [7:0] rowR_416;
wire [7:0] rowR_417;
wire [7:0] rowR_418;
wire [7:0] rowR_419;
wire [7:0] rowR_420;
wire [7:0] rowR_421;
wire [7:0] rowR_422;
wire [7:0] rowR_423;
wire [7:0] rowR_424;
wire [7:0] rowR_425;
wire [7:0] rowR_426;
wire [7:0] rowR_427;
wire [7:0] rowR_428;
wire [7:0] rowR_429;
wire [7:0] rowR_430;
wire [7:0] rowR_431;
wire [7:0] rowR_432;
wire [7:0] rowR_433;
wire [7:0] rowR_434;
wire [7:0] rowR_435;
wire [7:0] rowR_436;
wire [7:0] rowR_437;
wire [7:0] rowR_438;
wire [7:0] rowR_439;
wire [7:0] rowR_440;
wire [7:0] rowR_441;
wire [7:0] rowR_442;
wire [7:0] rowR_443;
wire [7:0] rowR_444;
wire [7:0] rowR_445;
wire [7:0] rowR_446;
wire [7:0] rowR_447;
wire [7:0] rowR_448;
wire [7:0] rowR_449;
wire [7:0] rowR_450;
wire [7:0] rowR_451;
wire [7:0] rowR_452;
wire [7:0] rowR_453;
wire [7:0] rowR_454;
wire [7:0] rowR_455;
wire [7:0] rowR_456;
wire [7:0] rowR_457;
wire [7:0] rowR_458;
wire [7:0] rowR_459;
wire [7:0] rowR_460;
wire [7:0] rowR_461;
wire [7:0] rowR_462;
wire [7:0] rowR_463;
wire [7:0] rowR_464;
wire [7:0] rowR_465;
wire [7:0] rowR_466;
wire [7:0] rowR_467;
wire [7:0] rowR_468;
wire [7:0] rowR_469;
wire [7:0] rowR_470;
wire [7:0] rowR_471;
wire [7:0] rowR_472;
wire [7:0] rowR_473;
wire [7:0] rowR_474;
wire [7:0] rowR_475;
wire [7:0] rowR_476;
wire [7:0] rowR_477;
wire [7:0] rowR_478;
wire [7:0] rowR_479;
wire [7:0] rowR_480;
wire [7:0] rowR_481;
wire [7:0] rowR_482;
wire [7:0] rowR_483;
wire [7:0] rowR_484;
wire [7:0] rowR_485;
wire [7:0] rowR_486;
wire [7:0] rowR_487;
wire [7:0] rowR_488;
wire [7:0] rowR_489;
wire [7:0] rowR_490;
wire [7:0] rowR_491;
wire [7:0] rowR_492;
wire [7:0] rowR_493;
wire [7:0] rowR_494;
wire [7:0] rowR_495;
wire [7:0] rowR_496;
wire [7:0] rowR_497;
wire [7:0] rowR_498;
wire [7:0] rowR_499;
wire [7:0] rowR_500;
wire [7:0] rowR_501;
wire [7:0] rowR_502;
wire [7:0] rowR_503;
wire [7:0] rowR_504;
wire [7:0] rowR_505;
wire [7:0] rowR_506;
wire [7:0] rowR_507;
wire [7:0] rowR_508;
wire [7:0] rowR_509;
wire [7:0] rowR_510;
wire [7:0] rowR_511;
wire [7:0] rowR_512;
wire [7:0] rowR_513;
wire [7:0] rowR_514;
wire [7:0] rowR_515;
wire [7:0] rowR_516;
wire [7:0] rowR_517;
wire [7:0] rowR_518;
wire [7:0] rowR_519;
wire [7:0] rowR_520;
wire [7:0] rowR_521;
wire [7:0] rowR_522;
wire [7:0] rowR_523;
wire [7:0] rowR_524;
wire [7:0] rowR_525;
wire [7:0] rowR_526;
wire [7:0] rowR_527;
wire [7:0] rowR_528;
wire [7:0] rowR_529;
wire [7:0] rowR_530;
wire [7:0] rowR_531;
wire [7:0] rowR_532;
wire [7:0] rowR_533;
wire [7:0] rowR_534;
wire [7:0] rowR_535;
wire [7:0] rowR_536;
wire [7:0] rowR_537;
wire [7:0] rowR_538;
wire [7:0] rowR_539;
wire [7:0] rowR_540;
wire [7:0] rowR_541;
wire [7:0] rowR_542;
wire [7:0] rowR_543;
wire [7:0] rowR_544;
wire [7:0] rowR_545;
wire [7:0] rowR_546;
wire [7:0] rowR_547;
wire [7:0] rowR_548;
wire [7:0] rowR_549;
wire [7:0] rowR_550;
wire [7:0] rowR_551;
wire [7:0] rowR_552;
wire [7:0] rowR_553;
wire [7:0] rowR_554;
wire [7:0] rowR_555;
wire [7:0] rowR_556;
wire [7:0] rowR_557;
wire [7:0] rowR_558;
wire [7:0] rowR_559;
wire [7:0] rowR_560;
wire [7:0] rowR_561;
wire [7:0] rowR_562;
wire [7:0] rowR_563;
wire [7:0] rowR_564;
wire [7:0] rowR_565;
wire [7:0] rowR_566;
wire [7:0] rowR_567;
wire [7:0] rowR_568;
wire [7:0] rowR_569;
wire [7:0] rowR_570;
wire [7:0] rowR_571;
wire [7:0] rowR_572;
wire [7:0] rowR_573;
wire [7:0] rowR_574;
wire [7:0] rowR_575;
wire [7:0] rowR_576;
wire [7:0] rowR_577;
wire [7:0] rowR_578;
wire [7:0] rowR_579;
wire [7:0] rowR_580;
wire [7:0] rowR_581;
wire [7:0] rowR_582;
wire [7:0] rowR_583;
wire [7:0] rowR_584;
wire [7:0] rowR_585;
wire [7:0] rowR_586;
wire [7:0] rowR_587;
wire [7:0] rowR_588;
wire [7:0] rowR_589;
wire [7:0] rowR_590;
wire [7:0] rowR_591;
wire [7:0] rowR_592;
wire [7:0] rowR_593;
wire [7:0] rowR_594;
wire [7:0] rowR_595;
wire [7:0] rowR_596;
wire [7:0] rowR_597;
wire [7:0] rowR_598;
wire [7:0] rowR_599;
wire [7:0] rowR_600;
wire [7:0] rowR_601;
wire [7:0] rowR_602;
wire [7:0] rowR_603;
wire [7:0] rowR_604;
wire [7:0] rowR_605;
wire [7:0] rowR_606;
wire [7:0] rowR_607;
wire [7:0] rowR_608;
wire [7:0] rowR_609;
wire [7:0] rowR_610;
wire [7:0] rowR_611;
wire [7:0] rowR_612;
wire [7:0] rowR_613;
wire [7:0] rowR_614;
wire [7:0] rowR_615;
wire [7:0] rowR_616;
wire [7:0] rowR_617;
wire [7:0] rowR_618;
wire [7:0] rowR_619;
wire [7:0] rowR_620;
wire [7:0] rowR_621;
wire [7:0] rowR_622;
wire [7:0] rowR_623;
wire [7:0] rowR_624;
wire [7:0] rowR_625;
wire [7:0] rowR_626;
wire [7:0] rowR_627;
wire [7:0] rowR_628;
wire [7:0] rowR_629;
wire [7:0] rowR_630;
wire [7:0] rowR_631;
wire [7:0] rowR_632;
wire [7:0] rowR_633;
wire [7:0] rowR_634;
wire [7:0] rowR_635;
wire [7:0] rowR_636;
wire [7:0] rowR_637;
wire [7:0] rowR_638;
wire [7:0] rowR_639;

wire [7:0] rowD_0;
wire [7:0] rowD_1;
wire [7:0] rowD_2;
wire [7:0] rowD_3;
wire [7:0] rowD_4;
wire [7:0] rowD_5;
wire [7:0] rowD_6;
wire [7:0] rowD_7;
wire [7:0] rowD_8;
wire [7:0] rowD_9;
wire [7:0] rowD_10;
wire [7:0] rowD_11;
wire [7:0] rowD_12;
wire [7:0] rowD_13;
wire [7:0] rowD_14;
wire [7:0] rowD_15;
wire [7:0] rowD_16;
wire [7:0] rowD_17;
wire [7:0] rowD_18;
wire [7:0] rowD_19;
wire [7:0] rowD_20;
wire [7:0] rowD_21;
wire [7:0] rowD_22;
wire [7:0] rowD_23;
wire [7:0] rowD_24;
wire [7:0] rowD_25;
wire [7:0] rowD_26;
wire [7:0] rowD_27;
wire [7:0] rowD_28;
wire [7:0] rowD_29;
wire [7:0] rowD_30;
wire [7:0] rowD_31;
wire [7:0] rowD_32;
wire [7:0] rowD_33;
wire [7:0] rowD_34;
wire [7:0] rowD_35;
wire [7:0] rowD_36;
wire [7:0] rowD_37;
wire [7:0] rowD_38;
wire [7:0] rowD_39;
wire [7:0] rowD_40;
wire [7:0] rowD_41;
wire [7:0] rowD_42;
wire [7:0] rowD_43;
wire [7:0] rowD_44;
wire [7:0] rowD_45;
wire [7:0] rowD_46;
wire [7:0] rowD_47;
wire [7:0] rowD_48;
wire [7:0] rowD_49;
wire [7:0] rowD_50;
wire [7:0] rowD_51;
wire [7:0] rowD_52;
wire [7:0] rowD_53;
wire [7:0] rowD_54;
wire [7:0] rowD_55;
wire [7:0] rowD_56;
wire [7:0] rowD_57;
wire [7:0] rowD_58;
wire [7:0] rowD_59;
wire [7:0] rowD_60;
wire [7:0] rowD_61;
wire [7:0] rowD_62;
wire [7:0] rowD_63;
wire [7:0] rowD_64;
wire [7:0] rowD_65;
wire [7:0] rowD_66;
wire [7:0] rowD_67;
wire [7:0] rowD_68;
wire [7:0] rowD_69;
wire [7:0] rowD_70;
wire [7:0] rowD_71;
wire [7:0] rowD_72;
wire [7:0] rowD_73;
wire [7:0] rowD_74;
wire [7:0] rowD_75;
wire [7:0] rowD_76;
wire [7:0] rowD_77;
wire [7:0] rowD_78;
wire [7:0] rowD_79;
wire [7:0] rowD_80;
wire [7:0] rowD_81;
wire [7:0] rowD_82;
wire [7:0] rowD_83;
wire [7:0] rowD_84;
wire [7:0] rowD_85;
wire [7:0] rowD_86;
wire [7:0] rowD_87;
wire [7:0] rowD_88;
wire [7:0] rowD_89;
wire [7:0] rowD_90;
wire [7:0] rowD_91;
wire [7:0] rowD_92;
wire [7:0] rowD_93;
wire [7:0] rowD_94;
wire [7:0] rowD_95;
wire [7:0] rowD_96;
wire [7:0] rowD_97;
wire [7:0] rowD_98;
wire [7:0] rowD_99;
wire [7:0] rowD_100;
wire [7:0] rowD_101;
wire [7:0] rowD_102;
wire [7:0] rowD_103;
wire [7:0] rowD_104;
wire [7:0] rowD_105;
wire [7:0] rowD_106;
wire [7:0] rowD_107;
wire [7:0] rowD_108;
wire [7:0] rowD_109;
wire [7:0] rowD_110;
wire [7:0] rowD_111;
wire [7:0] rowD_112;
wire [7:0] rowD_113;
wire [7:0] rowD_114;
wire [7:0] rowD_115;
wire [7:0] rowD_116;
wire [7:0] rowD_117;
wire [7:0] rowD_118;
wire [7:0] rowD_119;
wire [7:0] rowD_120;
wire [7:0] rowD_121;
wire [7:0] rowD_122;
wire [7:0] rowD_123;
wire [7:0] rowD_124;
wire [7:0] rowD_125;
wire [7:0] rowD_126;
wire [7:0] rowD_127;
wire [7:0] rowD_128;
wire [7:0] rowD_129;
wire [7:0] rowD_130;
wire [7:0] rowD_131;
wire [7:0] rowD_132;
wire [7:0] rowD_133;
wire [7:0] rowD_134;
wire [7:0] rowD_135;
wire [7:0] rowD_136;
wire [7:0] rowD_137;
wire [7:0] rowD_138;
wire [7:0] rowD_139;
wire [7:0] rowD_140;
wire [7:0] rowD_141;
wire [7:0] rowD_142;
wire [7:0] rowD_143;
wire [7:0] rowD_144;
wire [7:0] rowD_145;
wire [7:0] rowD_146;
wire [7:0] rowD_147;
wire [7:0] rowD_148;
wire [7:0] rowD_149;
wire [7:0] rowD_150;
wire [7:0] rowD_151;
wire [7:0] rowD_152;
wire [7:0] rowD_153;
wire [7:0] rowD_154;
wire [7:0] rowD_155;
wire [7:0] rowD_156;
wire [7:0] rowD_157;
wire [7:0] rowD_158;
wire [7:0] rowD_159;
wire [7:0] rowD_160;
wire [7:0] rowD_161;
wire [7:0] rowD_162;
wire [7:0] rowD_163;
wire [7:0] rowD_164;
wire [7:0] rowD_165;
wire [7:0] rowD_166;
wire [7:0] rowD_167;
wire [7:0] rowD_168;
wire [7:0] rowD_169;
wire [7:0] rowD_170;
wire [7:0] rowD_171;
wire [7:0] rowD_172;
wire [7:0] rowD_173;
wire [7:0] rowD_174;
wire [7:0] rowD_175;
wire [7:0] rowD_176;
wire [7:0] rowD_177;
wire [7:0] rowD_178;
wire [7:0] rowD_179;
wire [7:0] rowD_180;
wire [7:0] rowD_181;
wire [7:0] rowD_182;
wire [7:0] rowD_183;
wire [7:0] rowD_184;
wire [7:0] rowD_185;
wire [7:0] rowD_186;
wire [7:0] rowD_187;
wire [7:0] rowD_188;
wire [7:0] rowD_189;
wire [7:0] rowD_190;
wire [7:0] rowD_191;
wire [7:0] rowD_192;
wire [7:0] rowD_193;
wire [7:0] rowD_194;
wire [7:0] rowD_195;
wire [7:0] rowD_196;
wire [7:0] rowD_197;
wire [7:0] rowD_198;
wire [7:0] rowD_199;
wire [7:0] rowD_200;
wire [7:0] rowD_201;
wire [7:0] rowD_202;
wire [7:0] rowD_203;
wire [7:0] rowD_204;
wire [7:0] rowD_205;
wire [7:0] rowD_206;
wire [7:0] rowD_207;
wire [7:0] rowD_208;
wire [7:0] rowD_209;
wire [7:0] rowD_210;
wire [7:0] rowD_211;
wire [7:0] rowD_212;
wire [7:0] rowD_213;
wire [7:0] rowD_214;
wire [7:0] rowD_215;
wire [7:0] rowD_216;
wire [7:0] rowD_217;
wire [7:0] rowD_218;
wire [7:0] rowD_219;
wire [7:0] rowD_220;
wire [7:0] rowD_221;
wire [7:0] rowD_222;
wire [7:0] rowD_223;
wire [7:0] rowD_224;
wire [7:0] rowD_225;
wire [7:0] rowD_226;
wire [7:0] rowD_227;
wire [7:0] rowD_228;
wire [7:0] rowD_229;
wire [7:0] rowD_230;
wire [7:0] rowD_231;
wire [7:0] rowD_232;
wire [7:0] rowD_233;
wire [7:0] rowD_234;
wire [7:0] rowD_235;
wire [7:0] rowD_236;
wire [7:0] rowD_237;
wire [7:0] rowD_238;
wire [7:0] rowD_239;
wire [7:0] rowD_240;
wire [7:0] rowD_241;
wire [7:0] rowD_242;
wire [7:0] rowD_243;
wire [7:0] rowD_244;
wire [7:0] rowD_245;
wire [7:0] rowD_246;
wire [7:0] rowD_247;
wire [7:0] rowD_248;
wire [7:0] rowD_249;
wire [7:0] rowD_250;
wire [7:0] rowD_251;
wire [7:0] rowD_252;
wire [7:0] rowD_253;
wire [7:0] rowD_254;
wire [7:0] rowD_255;
wire [7:0] rowD_256;
wire [7:0] rowD_257;
wire [7:0] rowD_258;
wire [7:0] rowD_259;
wire [7:0] rowD_260;
wire [7:0] rowD_261;
wire [7:0] rowD_262;
wire [7:0] rowD_263;
wire [7:0] rowD_264;
wire [7:0] rowD_265;
wire [7:0] rowD_266;
wire [7:0] rowD_267;
wire [7:0] rowD_268;
wire [7:0] rowD_269;
wire [7:0] rowD_270;
wire [7:0] rowD_271;
wire [7:0] rowD_272;
wire [7:0] rowD_273;
wire [7:0] rowD_274;
wire [7:0] rowD_275;
wire [7:0] rowD_276;
wire [7:0] rowD_277;
wire [7:0] rowD_278;
wire [7:0] rowD_279;
wire [7:0] rowD_280;
wire [7:0] rowD_281;
wire [7:0] rowD_282;
wire [7:0] rowD_283;
wire [7:0] rowD_284;
wire [7:0] rowD_285;
wire [7:0] rowD_286;
wire [7:0] rowD_287;
wire [7:0] rowD_288;
wire [7:0] rowD_289;
wire [7:0] rowD_290;
wire [7:0] rowD_291;
wire [7:0] rowD_292;
wire [7:0] rowD_293;
wire [7:0] rowD_294;
wire [7:0] rowD_295;
wire [7:0] rowD_296;
wire [7:0] rowD_297;
wire [7:0] rowD_298;
wire [7:0] rowD_299;
wire [7:0] rowD_300;
wire [7:0] rowD_301;
wire [7:0] rowD_302;
wire [7:0] rowD_303;
wire [7:0] rowD_304;
wire [7:0] rowD_305;
wire [7:0] rowD_306;
wire [7:0] rowD_307;
wire [7:0] rowD_308;
wire [7:0] rowD_309;
wire [7:0] rowD_310;
wire [7:0] rowD_311;
wire [7:0] rowD_312;
wire [7:0] rowD_313;
wire [7:0] rowD_314;
wire [7:0] rowD_315;
wire [7:0] rowD_316;
wire [7:0] rowD_317;
wire [7:0] rowD_318;
wire [7:0] rowD_319;
wire [7:0] rowD_320;
wire [7:0] rowD_321;
wire [7:0] rowD_322;
wire [7:0] rowD_323;
wire [7:0] rowD_324;
wire [7:0] rowD_325;
wire [7:0] rowD_326;
wire [7:0] rowD_327;
wire [7:0] rowD_328;
wire [7:0] rowD_329;
wire [7:0] rowD_330;
wire [7:0] rowD_331;
wire [7:0] rowD_332;
wire [7:0] rowD_333;
wire [7:0] rowD_334;
wire [7:0] rowD_335;
wire [7:0] rowD_336;
wire [7:0] rowD_337;
wire [7:0] rowD_338;
wire [7:0] rowD_339;
wire [7:0] rowD_340;
wire [7:0] rowD_341;
wire [7:0] rowD_342;
wire [7:0] rowD_343;
wire [7:0] rowD_344;
wire [7:0] rowD_345;
wire [7:0] rowD_346;
wire [7:0] rowD_347;
wire [7:0] rowD_348;
wire [7:0] rowD_349;
wire [7:0] rowD_350;
wire [7:0] rowD_351;
wire [7:0] rowD_352;
wire [7:0] rowD_353;
wire [7:0] rowD_354;
wire [7:0] rowD_355;
wire [7:0] rowD_356;
wire [7:0] rowD_357;
wire [7:0] rowD_358;
wire [7:0] rowD_359;
wire [7:0] rowD_360;
wire [7:0] rowD_361;
wire [7:0] rowD_362;
wire [7:0] rowD_363;
wire [7:0] rowD_364;
wire [7:0] rowD_365;
wire [7:0] rowD_366;
wire [7:0] rowD_367;
wire [7:0] rowD_368;
wire [7:0] rowD_369;
wire [7:0] rowD_370;
wire [7:0] rowD_371;
wire [7:0] rowD_372;
wire [7:0] rowD_373;
wire [7:0] rowD_374;
wire [7:0] rowD_375;
wire [7:0] rowD_376;
wire [7:0] rowD_377;
wire [7:0] rowD_378;
wire [7:0] rowD_379;
wire [7:0] rowD_380;
wire [7:0] rowD_381;
wire [7:0] rowD_382;
wire [7:0] rowD_383;
wire [7:0] rowD_384;
wire [7:0] rowD_385;
wire [7:0] rowD_386;
wire [7:0] rowD_387;
wire [7:0] rowD_388;
wire [7:0] rowD_389;
wire [7:0] rowD_390;
wire [7:0] rowD_391;
wire [7:0] rowD_392;
wire [7:0] rowD_393;
wire [7:0] rowD_394;
wire [7:0] rowD_395;
wire [7:0] rowD_396;
wire [7:0] rowD_397;
wire [7:0] rowD_398;
wire [7:0] rowD_399;
wire [7:0] rowD_400;
wire [7:0] rowD_401;
wire [7:0] rowD_402;
wire [7:0] rowD_403;
wire [7:0] rowD_404;
wire [7:0] rowD_405;
wire [7:0] rowD_406;
wire [7:0] rowD_407;
wire [7:0] rowD_408;
wire [7:0] rowD_409;
wire [7:0] rowD_410;
wire [7:0] rowD_411;
wire [7:0] rowD_412;
wire [7:0] rowD_413;
wire [7:0] rowD_414;
wire [7:0] rowD_415;
wire [7:0] rowD_416;
wire [7:0] rowD_417;
wire [7:0] rowD_418;
wire [7:0] rowD_419;
wire [7:0] rowD_420;
wire [7:0] rowD_421;
wire [7:0] rowD_422;
wire [7:0] rowD_423;
wire [7:0] rowD_424;
wire [7:0] rowD_425;
wire [7:0] rowD_426;
wire [7:0] rowD_427;
wire [7:0] rowD_428;
wire [7:0] rowD_429;
wire [7:0] rowD_430;
wire [7:0] rowD_431;
wire [7:0] rowD_432;
wire [7:0] rowD_433;
wire [7:0] rowD_434;
wire [7:0] rowD_435;
wire [7:0] rowD_436;
wire [7:0] rowD_437;
wire [7:0] rowD_438;
wire [7:0] rowD_439;
wire [7:0] rowD_440;
wire [7:0] rowD_441;
wire [7:0] rowD_442;
wire [7:0] rowD_443;
wire [7:0] rowD_444;
wire [7:0] rowD_445;
wire [7:0] rowD_446;
wire [7:0] rowD_447;
wire [7:0] rowD_448;
wire [7:0] rowD_449;
wire [7:0] rowD_450;
wire [7:0] rowD_451;
wire [7:0] rowD_452;
wire [7:0] rowD_453;
wire [7:0] rowD_454;
wire [7:0] rowD_455;
wire [7:0] rowD_456;
wire [7:0] rowD_457;
wire [7:0] rowD_458;
wire [7:0] rowD_459;
wire [7:0] rowD_460;
wire [7:0] rowD_461;
wire [7:0] rowD_462;
wire [7:0] rowD_463;
wire [7:0] rowD_464;
wire [7:0] rowD_465;
wire [7:0] rowD_466;
wire [7:0] rowD_467;
wire [7:0] rowD_468;
wire [7:0] rowD_469;
wire [7:0] rowD_470;
wire [7:0] rowD_471;
wire [7:0] rowD_472;
wire [7:0] rowD_473;
wire [7:0] rowD_474;
wire [7:0] rowD_475;
wire [7:0] rowD_476;
wire [7:0] rowD_477;
wire [7:0] rowD_478;
wire [7:0] rowD_479;
wire [7:0] rowD_480;
wire [7:0] rowD_481;
wire [7:0] rowD_482;
wire [7:0] rowD_483;
wire [7:0] rowD_484;
wire [7:0] rowD_485;
wire [7:0] rowD_486;
wire [7:0] rowD_487;
wire [7:0] rowD_488;
wire [7:0] rowD_489;
wire [7:0] rowD_490;
wire [7:0] rowD_491;
wire [7:0] rowD_492;
wire [7:0] rowD_493;
wire [7:0] rowD_494;
wire [7:0] rowD_495;
wire [7:0] rowD_496;
wire [7:0] rowD_497;
wire [7:0] rowD_498;
wire [7:0] rowD_499;
wire [7:0] rowD_500;
wire [7:0] rowD_501;
wire [7:0] rowD_502;
wire [7:0] rowD_503;
wire [7:0] rowD_504;
wire [7:0] rowD_505;
wire [7:0] rowD_506;
wire [7:0] rowD_507;
wire [7:0] rowD_508;
wire [7:0] rowD_509;
wire [7:0] rowD_510;
wire [7:0] rowD_511;
wire [7:0] rowD_512;
wire [7:0] rowD_513;
wire [7:0] rowD_514;
wire [7:0] rowD_515;
wire [7:0] rowD_516;
wire [7:0] rowD_517;
wire [7:0] rowD_518;
wire [7:0] rowD_519;
wire [7:0] rowD_520;
wire [7:0] rowD_521;
wire [7:0] rowD_522;
wire [7:0] rowD_523;
wire [7:0] rowD_524;
wire [7:0] rowD_525;
wire [7:0] rowD_526;
wire [7:0] rowD_527;
wire [7:0] rowD_528;
wire [7:0] rowD_529;
wire [7:0] rowD_530;
wire [7:0] rowD_531;
wire [7:0] rowD_532;
wire [7:0] rowD_533;
wire [7:0] rowD_534;
wire [7:0] rowD_535;
wire [7:0] rowD_536;
wire [7:0] rowD_537;
wire [7:0] rowD_538;
wire [7:0] rowD_539;
wire [7:0] rowD_540;
wire [7:0] rowD_541;
wire [7:0] rowD_542;
wire [7:0] rowD_543;
wire [7:0] rowD_544;
wire [7:0] rowD_545;
wire [7:0] rowD_546;
wire [7:0] rowD_547;
wire [7:0] rowD_548;
wire [7:0] rowD_549;
wire [7:0] rowD_550;
wire [7:0] rowD_551;
wire [7:0] rowD_552;
wire [7:0] rowD_553;
wire [7:0] rowD_554;
wire [7:0] rowD_555;
wire [7:0] rowD_556;
wire [7:0] rowD_557;
wire [7:0] rowD_558;
wire [7:0] rowD_559;
wire [7:0] rowD_560;
wire [7:0] rowD_561;
wire [7:0] rowD_562;
wire [7:0] rowD_563;
wire [7:0] rowD_564;
wire [7:0] rowD_565;
wire [7:0] rowD_566;
wire [7:0] rowD_567;
wire [7:0] rowD_568;
wire [7:0] rowD_569;
wire [7:0] rowD_570;
wire [7:0] rowD_571;
wire [7:0] rowD_572;
wire [7:0] rowD_573;
wire [7:0] rowD_574;
wire [7:0] rowD_575;
wire [7:0] rowD_576;
wire [7:0] rowD_577;
wire [7:0] rowD_578;
wire [7:0] rowD_579;
wire [7:0] rowD_580;
wire [7:0] rowD_581;
wire [7:0] rowD_582;
wire [7:0] rowD_583;
wire [7:0] rowD_584;
wire [7:0] rowD_585;
wire [7:0] rowD_586;
wire [7:0] rowD_587;
wire [7:0] rowD_588;
wire [7:0] rowD_589;
wire [7:0] rowD_590;
wire [7:0] rowD_591;
wire [7:0] rowD_592;
wire [7:0] rowD_593;
wire [7:0] rowD_594;
wire [7:0] rowD_595;
wire [7:0] rowD_596;
wire [7:0] rowD_597;
wire [7:0] rowD_598;
wire [7:0] rowD_599;
wire [7:0] rowD_600;
wire [7:0] rowD_601;
wire [7:0] rowD_602;
wire [7:0] rowD_603;
wire [7:0] rowD_604;
wire [7:0] rowD_605;
wire [7:0] rowD_606;
wire [7:0] rowD_607;
wire [7:0] rowD_608;
wire [7:0] rowD_609;
wire [7:0] rowD_610;
wire [7:0] rowD_611;
wire [7:0] rowD_612;
wire [7:0] rowD_613;
wire [7:0] rowD_614;
wire [7:0] rowD_615;
wire [7:0] rowD_616;
wire [7:0] rowD_617;
wire [7:0] rowD_618;
wire [7:0] rowD_619;
wire [7:0] rowD_620;
wire [7:0] rowD_621;
wire [7:0] rowD_622;
wire [7:0] rowD_623;
wire [7:0] rowD_624;
wire [7:0] rowD_625;
wire [7:0] rowD_626;
wire [7:0] rowD_627;
wire [7:0] rowD_628;
wire [7:0] rowD_629;
wire [7:0] rowD_630;
wire [7:0] rowD_631;
wire [7:0] rowD_632;
wire [7:0] rowD_633;
wire [7:0] rowD_634;
wire [7:0] rowD_635;
wire [7:0] rowD_636;
wire [7:0] rowD_637;
wire [7:0] rowD_638;
wire [7:0] rowD_639;

wire enS2P1;
wire enS2P2;
wire enC;
wire enP2S;
wire enout;

wire ce_out1;
wire ce_out2;
wire ce_out3;
wire ce_out4;

Serial_to_Parallel_fixpt sp1
           (clk,
           reset,
           clk_enable,
           pixelL_in,
           ce_out1,
           rowL_0,
           rowL_1,
           rowL_2,
           rowL_3,
           rowL_4,
           rowL_5,
           rowL_6,
           rowL_7,
           rowL_8,
           rowL_9,
           rowL_10,
           rowL_11,
           rowL_12,
           rowL_13,
           rowL_14,
           rowL_15,
           rowL_16,
           rowL_17,
           rowL_18,
           rowL_19,
           rowL_20,
           rowL_21,
           rowL_22,
           rowL_23,
           rowL_24,
           rowL_25,
           rowL_26,
           rowL_27,
           rowL_28,
           rowL_29,
           rowL_30,
           rowL_31,
           rowL_32,
           rowL_33,
           rowL_34,
           rowL_35,
           rowL_36,
           rowL_37,
           rowL_38,
           rowL_39,
           rowL_40,
           rowL_41,
           rowL_42,
           rowL_43,
           rowL_44,
           rowL_45,
           rowL_46,
           rowL_47,
           rowL_48,
           rowL_49,
           rowL_50,
           rowL_51,
           rowL_52,
           rowL_53,
           rowL_54,
           rowL_55,
           rowL_56,
           rowL_57,
           rowL_58,
           rowL_59,
           rowL_60,
           rowL_61,
           rowL_62,
           rowL_63,
           rowL_64,
           rowL_65,
           rowL_66,
           rowL_67,
           rowL_68,
           rowL_69,
           rowL_70,
           rowL_71,
           rowL_72,
           rowL_73,
           rowL_74,
           rowL_75,
           rowL_76,
           rowL_77,
           rowL_78,
           rowL_79,
           rowL_80,
           rowL_81,
           rowL_82,
           rowL_83,
           rowL_84,
           rowL_85,
           rowL_86,
           rowL_87,
           rowL_88,
           rowL_89,
           rowL_90,
           rowL_91,
           rowL_92,
           rowL_93,
           rowL_94,
           rowL_95,
           rowL_96,
           rowL_97,
           rowL_98,
           rowL_99,
           rowL_100,
           rowL_101,
           rowL_102,
           rowL_103,
           rowL_104,
           rowL_105,
           rowL_106,
           rowL_107,
           rowL_108,
           rowL_109,
           rowL_110,
           rowL_111,
           rowL_112,
           rowL_113,
           rowL_114,
           rowL_115,
           rowL_116,
           rowL_117,
           rowL_118,
           rowL_119,
           rowL_120,
           rowL_121,
           rowL_122,
           rowL_123,
           rowL_124,
           rowL_125,
           rowL_126,
           rowL_127,
           rowL_128,
           rowL_129,
           rowL_130,
           rowL_131,
           rowL_132,
           rowL_133,
           rowL_134,
           rowL_135,
           rowL_136,
           rowL_137,
           rowL_138,
           rowL_139,
           rowL_140,
           rowL_141,
           rowL_142,
           rowL_143,
           rowL_144,
           rowL_145,
           rowL_146,
           rowL_147,
           rowL_148,
           rowL_149,
           rowL_150,
           rowL_151,
           rowL_152,
           rowL_153,
           rowL_154,
           rowL_155,
           rowL_156,
           rowL_157,
           rowL_158,
           rowL_159,
           rowL_160,
           rowL_161,
           rowL_162,
           rowL_163,
           rowL_164,
           rowL_165,
           rowL_166,
           rowL_167,
           rowL_168,
           rowL_169,
           rowL_170,
           rowL_171,
           rowL_172,
           rowL_173,
           rowL_174,
           rowL_175,
           rowL_176,
           rowL_177,
           rowL_178,
           rowL_179,
           rowL_180,
           rowL_181,
           rowL_182,
           rowL_183,
           rowL_184,
           rowL_185,
           rowL_186,
           rowL_187,
           rowL_188,
           rowL_189,
           rowL_190,
           rowL_191,
           rowL_192,
           rowL_193,
           rowL_194,
           rowL_195,
           rowL_196,
           rowL_197,
           rowL_198,
           rowL_199,
           rowL_200,
           rowL_201,
           rowL_202,
           rowL_203,
           rowL_204,
           rowL_205,
           rowL_206,
           rowL_207,
           rowL_208,
           rowL_209,
           rowL_210,
           rowL_211,
           rowL_212,
           rowL_213,
           rowL_214,
           rowL_215,
           rowL_216,
           rowL_217,
           rowL_218,
           rowL_219,
           rowL_220,
           rowL_221,
           rowL_222,
           rowL_223,
           rowL_224,
           rowL_225,
           rowL_226,
           rowL_227,
           rowL_228,
           rowL_229,
           rowL_230,
           rowL_231,
           rowL_232,
           rowL_233,
           rowL_234,
           rowL_235,
           rowL_236,
           rowL_237,
           rowL_238,
           rowL_239,
           rowL_240,
           rowL_241,
           rowL_242,
           rowL_243,
           rowL_244,
           rowL_245,
           rowL_246,
           rowL_247,
           rowL_248,
           rowL_249,
           rowL_250,
           rowL_251,
           rowL_252,
           rowL_253,
           rowL_254,
           rowL_255,
           rowL_256,
           rowL_257,
           rowL_258,
           rowL_259,
           rowL_260,
           rowL_261,
           rowL_262,
           rowL_263,
           rowL_264,
           rowL_265,
           rowL_266,
           rowL_267,
           rowL_268,
           rowL_269,
           rowL_270,
           rowL_271,
           rowL_272,
           rowL_273,
           rowL_274,
           rowL_275,
           rowL_276,
           rowL_277,
           rowL_278,
           rowL_279,
           rowL_280,
           rowL_281,
           rowL_282,
           rowL_283,
           rowL_284,
           rowL_285,
           rowL_286,
           rowL_287,
           rowL_288,
           rowL_289,
           rowL_290,
           rowL_291,
           rowL_292,
           rowL_293,
           rowL_294,
           rowL_295,
           rowL_296,
           rowL_297,
           rowL_298,
           rowL_299,
           rowL_300,
           rowL_301,
           rowL_302,
           rowL_303,
           rowL_304,
           rowL_305,
           rowL_306,
           rowL_307,
           rowL_308,
           rowL_309,
           rowL_310,
           rowL_311,
           rowL_312,
           rowL_313,
           rowL_314,
           rowL_315,
           rowL_316,
           rowL_317,
           rowL_318,
           rowL_319,
           rowL_320,
           rowL_321,
           rowL_322,
           rowL_323,
           rowL_324,
           rowL_325,
           rowL_326,
           rowL_327,
           rowL_328,
           rowL_329,
           rowL_330,
           rowL_331,
           rowL_332,
           rowL_333,
           rowL_334,
           rowL_335,
           rowL_336,
           rowL_337,
           rowL_338,
           rowL_339,
           rowL_340,
           rowL_341,
           rowL_342,
           rowL_343,
           rowL_344,
           rowL_345,
           rowL_346,
           rowL_347,
           rowL_348,
           rowL_349,
           rowL_350,
           rowL_351,
           rowL_352,
           rowL_353,
           rowL_354,
           rowL_355,
           rowL_356,
           rowL_357,
           rowL_358,
           rowL_359,
           rowL_360,
           rowL_361,
           rowL_362,
           rowL_363,
           rowL_364,
           rowL_365,
           rowL_366,
           rowL_367,
           rowL_368,
           rowL_369,
           rowL_370,
           rowL_371,
           rowL_372,
           rowL_373,
           rowL_374,
           rowL_375,
           rowL_376,
           rowL_377,
           rowL_378,
           rowL_379,
           rowL_380,
           rowL_381,
           rowL_382,
           rowL_383,
           rowL_384,
           rowL_385,
           rowL_386,
           rowL_387,
           rowL_388,
           rowL_389,
           rowL_390,
           rowL_391,
           rowL_392,
           rowL_393,
           rowL_394,
           rowL_395,
           rowL_396,
           rowL_397,
           rowL_398,
           rowL_399,
           rowL_400,
           rowL_401,
           rowL_402,
           rowL_403,
           rowL_404,
           rowL_405,
           rowL_406,
           rowL_407,
           rowL_408,
           rowL_409,
           rowL_410,
           rowL_411,
           rowL_412,
           rowL_413,
           rowL_414,
           rowL_415,
           rowL_416,
           rowL_417,
           rowL_418,
           rowL_419,
           rowL_420,
           rowL_421,
           rowL_422,
           rowL_423,
           rowL_424,
           rowL_425,
           rowL_426,
           rowL_427,
           rowL_428,
           rowL_429,
           rowL_430,
           rowL_431,
           rowL_432,
           rowL_433,
           rowL_434,
           rowL_435,
           rowL_436,
           rowL_437,
           rowL_438,
           rowL_439,
           rowL_440,
           rowL_441,
           rowL_442,
           rowL_443,
           rowL_444,
           rowL_445,
           rowL_446,
           rowL_447,
           rowL_448,
           rowL_449,
           rowL_450,
           rowL_451,
           rowL_452,
           rowL_453,
           rowL_454,
           rowL_455,
           rowL_456,
           rowL_457,
           rowL_458,
           rowL_459,
           rowL_460,
           rowL_461,
           rowL_462,
           rowL_463,
           rowL_464,
           rowL_465,
           rowL_466,
           rowL_467,
           rowL_468,
           rowL_469,
           rowL_470,
           rowL_471,
           rowL_472,
           rowL_473,
           rowL_474,
           rowL_475,
           rowL_476,
           rowL_477,
           rowL_478,
           rowL_479,
           rowL_480,
           rowL_481,
           rowL_482,
           rowL_483,
           rowL_484,
           rowL_485,
           rowL_486,
           rowL_487,
           rowL_488,
           rowL_489,
           rowL_490,
           rowL_491,
           rowL_492,
           rowL_493,
           rowL_494,
           rowL_495,
           rowL_496,
           rowL_497,
           rowL_498,
           rowL_499,
           rowL_500,
           rowL_501,
           rowL_502,
           rowL_503,
           rowL_504,
           rowL_505,
           rowL_506,
           rowL_507,
           rowL_508,
           rowL_509,
           rowL_510,
           rowL_511,
           rowL_512,
           rowL_513,
           rowL_514,
           rowL_515,
           rowL_516,
           rowL_517,
           rowL_518,
           rowL_519,
           rowL_520,
           rowL_521,
           rowL_522,
           rowL_523,
           rowL_524,
           rowL_525,
           rowL_526,
           rowL_527,
           rowL_528,
           rowL_529,
           rowL_530,
           rowL_531,
           rowL_532,
           rowL_533,
           rowL_534,
           rowL_535,
           rowL_536,
           rowL_537,
           rowL_538,
           rowL_539,
           rowL_540,
           rowL_541,
           rowL_542,
           rowL_543,
           rowL_544,
           rowL_545,
           rowL_546,
           rowL_547,
           rowL_548,
           rowL_549,
           rowL_550,
           rowL_551,
           rowL_552,
           rowL_553,
           rowL_554,
           rowL_555,
           rowL_556,
           rowL_557,
           rowL_558,
           rowL_559,
           rowL_560,
           rowL_561,
           rowL_562,
           rowL_563,
           rowL_564,
           rowL_565,
           rowL_566,
           rowL_567,
           rowL_568,
           rowL_569,
           rowL_570,
           rowL_571,
           rowL_572,
           rowL_573,
           rowL_574,
           rowL_575,
           rowL_576,
           rowL_577,
           rowL_578,
           rowL_579,
           rowL_580,
           rowL_581,
           rowL_582,
           rowL_583,
           rowL_584,
           rowL_585,
           rowL_586,
           rowL_587,
           rowL_588,
           rowL_589,
           rowL_590,
           rowL_591,
           rowL_592,
           rowL_593,
           rowL_594,
           rowL_595,
           rowL_596,
           rowL_597,
           rowL_598,
           rowL_599,
           rowL_600,
           rowL_601,
           rowL_602,
           rowL_603,
           rowL_604,
           rowL_605,
           rowL_606,
           rowL_607,
           rowL_608,
           rowL_609,
           rowL_610,
           rowL_611,
           rowL_612,
           rowL_613,
           rowL_614,
           rowL_615,
           rowL_616,
           rowL_617,
           rowL_618,
           rowL_619,
           rowL_620,
           rowL_621,
           rowL_622,
           rowL_623,
           rowL_624,
           rowL_625,
           rowL_626,
           rowL_627,
           rowL_628,
           rowL_629,
           rowL_630,
           rowL_631,
           rowL_632,
           rowL_633,
           rowL_634,
           rowL_635,
           rowL_636,
           rowL_637,
           rowL_638,
           rowL_639,
           enS2P1
);

Serial_to_Parallel_fixpt sp2
           (clk,
           reset,
           clk_enable,
           pixelR_in,
           ce_out2,
           rowR_0,
           rowR_1,
           rowR_2,
           rowR_3,
           rowR_4,
           rowR_5,
           rowR_6,
           rowR_7,
           rowR_8,
           rowR_9,
           rowR_10,
           rowR_11,
           rowR_12,
           rowR_13,
           rowR_14,
           rowR_15,
           rowR_16,
           rowR_17,
           rowR_18,
           rowR_19,
           rowR_20,
           rowR_21,
           rowR_22,
           rowR_23,
           rowR_24,
           rowR_25,
           rowR_26,
           rowR_27,
           rowR_28,
           rowR_29,
           rowR_30,
           rowR_31,
           rowR_32,
           rowR_33,
           rowR_34,
           rowR_35,
           rowR_36,
           rowR_37,
           rowR_38,
           rowR_39,
           rowR_40,
           rowR_41,
           rowR_42,
           rowR_43,
           rowR_44,
           rowR_45,
           rowR_46,
           rowR_47,
           rowR_48,
           rowR_49,
           rowR_50,
           rowR_51,
           rowR_52,
           rowR_53,
           rowR_54,
           rowR_55,
           rowR_56,
           rowR_57,
           rowR_58,
           rowR_59,
           rowR_60,
           rowR_61,
           rowR_62,
           rowR_63,
           rowR_64,
           rowR_65,
           rowR_66,
           rowR_67,
           rowR_68,
           rowR_69,
           rowR_70,
           rowR_71,
           rowR_72,
           rowR_73,
           rowR_74,
           rowR_75,
           rowR_76,
           rowR_77,
           rowR_78,
           rowR_79,
           rowR_80,
           rowR_81,
           rowR_82,
           rowR_83,
           rowR_84,
           rowR_85,
           rowR_86,
           rowR_87,
           rowR_88,
           rowR_89,
           rowR_90,
           rowR_91,
           rowR_92,
           rowR_93,
           rowR_94,
           rowR_95,
           rowR_96,
           rowR_97,
           rowR_98,
           rowR_99,
           rowR_100,
           rowR_101,
           rowR_102,
           rowR_103,
           rowR_104,
           rowR_105,
           rowR_106,
           rowR_107,
           rowR_108,
           rowR_109,
           rowR_110,
           rowR_111,
           rowR_112,
           rowR_113,
           rowR_114,
           rowR_115,
           rowR_116,
           rowR_117,
           rowR_118,
           rowR_119,
           rowR_120,
           rowR_121,
           rowR_122,
           rowR_123,
           rowR_124,
           rowR_125,
           rowR_126,
           rowR_127,
           rowR_128,
           rowR_129,
           rowR_130,
           rowR_131,
           rowR_132,
           rowR_133,
           rowR_134,
           rowR_135,
           rowR_136,
           rowR_137,
           rowR_138,
           rowR_139,
           rowR_140,
           rowR_141,
           rowR_142,
           rowR_143,
           rowR_144,
           rowR_145,
           rowR_146,
           rowR_147,
           rowR_148,
           rowR_149,
           rowR_150,
           rowR_151,
           rowR_152,
           rowR_153,
           rowR_154,
           rowR_155,
           rowR_156,
           rowR_157,
           rowR_158,
           rowR_159,
           rowR_160,
           rowR_161,
           rowR_162,
           rowR_163,
           rowR_164,
           rowR_165,
           rowR_166,
           rowR_167,
           rowR_168,
           rowR_169,
           rowR_170,
           rowR_171,
           rowR_172,
           rowR_173,
           rowR_174,
           rowR_175,
           rowR_176,
           rowR_177,
           rowR_178,
           rowR_179,
           rowR_180,
           rowR_181,
           rowR_182,
           rowR_183,
           rowR_184,
           rowR_185,
           rowR_186,
           rowR_187,
           rowR_188,
           rowR_189,
           rowR_190,
           rowR_191,
           rowR_192,
           rowR_193,
           rowR_194,
           rowR_195,
           rowR_196,
           rowR_197,
           rowR_198,
           rowR_199,
           rowR_200,
           rowR_201,
           rowR_202,
           rowR_203,
           rowR_204,
           rowR_205,
           rowR_206,
           rowR_207,
           rowR_208,
           rowR_209,
           rowR_210,
           rowR_211,
           rowR_212,
           rowR_213,
           rowR_214,
           rowR_215,
           rowR_216,
           rowR_217,
           rowR_218,
           rowR_219,
           rowR_220,
           rowR_221,
           rowR_222,
           rowR_223,
           rowR_224,
           rowR_225,
           rowR_226,
           rowR_227,
           rowR_228,
           rowR_229,
           rowR_230,
           rowR_231,
           rowR_232,
           rowR_233,
           rowR_234,
           rowR_235,
           rowR_236,
           rowR_237,
           rowR_238,
           rowR_239,
           rowR_240,
           rowR_241,
           rowR_242,
           rowR_243,
           rowR_244,
           rowR_245,
           rowR_246,
           rowR_247,
           rowR_248,
           rowR_249,
           rowR_250,
           rowR_251,
           rowR_252,
           rowR_253,
           rowR_254,
           rowR_255,
           rowR_256,
           rowR_257,
           rowR_258,
           rowR_259,
           rowR_260,
           rowR_261,
           rowR_262,
           rowR_263,
           rowR_264,
           rowR_265,
           rowR_266,
           rowR_267,
           rowR_268,
           rowR_269,
           rowR_270,
           rowR_271,
           rowR_272,
           rowR_273,
           rowR_274,
           rowR_275,
           rowR_276,
           rowR_277,
           rowR_278,
           rowR_279,
           rowR_280,
           rowR_281,
           rowR_282,
           rowR_283,
           rowR_284,
           rowR_285,
           rowR_286,
           rowR_287,
           rowR_288,
           rowR_289,
           rowR_290,
           rowR_291,
           rowR_292,
           rowR_293,
           rowR_294,
           rowR_295,
           rowR_296,
           rowR_297,
           rowR_298,
           rowR_299,
           rowR_300,
           rowR_301,
           rowR_302,
           rowR_303,
           rowR_304,
           rowR_305,
           rowR_306,
           rowR_307,
           rowR_308,
           rowR_309,
           rowR_310,
           rowR_311,
           rowR_312,
           rowR_313,
           rowR_314,
           rowR_315,
           rowR_316,
           rowR_317,
           rowR_318,
           rowR_319,
           rowR_320,
           rowR_321,
           rowR_322,
           rowR_323,
           rowR_324,
           rowR_325,
           rowR_326,
           rowR_327,
           rowR_328,
           rowR_329,
           rowR_330,
           rowR_331,
           rowR_332,
           rowR_333,
           rowR_334,
           rowR_335,
           rowR_336,
           rowR_337,
           rowR_338,
           rowR_339,
           rowR_340,
           rowR_341,
           rowR_342,
           rowR_343,
           rowR_344,
           rowR_345,
           rowR_346,
           rowR_347,
           rowR_348,
           rowR_349,
           rowR_350,
           rowR_351,
           rowR_352,
           rowR_353,
           rowR_354,
           rowR_355,
           rowR_356,
           rowR_357,
           rowR_358,
           rowR_359,
           rowR_360,
           rowR_361,
           rowR_362,
           rowR_363,
           rowR_364,
           rowR_365,
           rowR_366,
           rowR_367,
           rowR_368,
           rowR_369,
           rowR_370,
           rowR_371,
           rowR_372,
           rowR_373,
           rowR_374,
           rowR_375,
           rowR_376,
           rowR_377,
           rowR_378,
           rowR_379,
           rowR_380,
           rowR_381,
           rowR_382,
           rowR_383,
           rowR_384,
           rowR_385,
           rowR_386,
           rowR_387,
           rowR_388,
           rowR_389,
           rowR_390,
           rowR_391,
           rowR_392,
           rowR_393,
           rowR_394,
           rowR_395,
           rowR_396,
           rowR_397,
           rowR_398,
           rowR_399,
           rowR_400,
           rowR_401,
           rowR_402,
           rowR_403,
           rowR_404,
           rowR_405,
           rowR_406,
           rowR_407,
           rowR_408,
           rowR_409,
           rowR_410,
           rowR_411,
           rowR_412,
           rowR_413,
           rowR_414,
           rowR_415,
           rowR_416,
           rowR_417,
           rowR_418,
           rowR_419,
           rowR_420,
           rowR_421,
           rowR_422,
           rowR_423,
           rowR_424,
           rowR_425,
           rowR_426,
           rowR_427,
           rowR_428,
           rowR_429,
           rowR_430,
           rowR_431,
           rowR_432,
           rowR_433,
           rowR_434,
           rowR_435,
           rowR_436,
           rowR_437,
           rowR_438,
           rowR_439,
           rowR_440,
           rowR_441,
           rowR_442,
           rowR_443,
           rowR_444,
           rowR_445,
           rowR_446,
           rowR_447,
           rowR_448,
           rowR_449,
           rowR_450,
           rowR_451,
           rowR_452,
           rowR_453,
           rowR_454,
           rowR_455,
           rowR_456,
           rowR_457,
           rowR_458,
           rowR_459,
           rowR_460,
           rowR_461,
           rowR_462,
           rowR_463,
           rowR_464,
           rowR_465,
           rowR_466,
           rowR_467,
           rowR_468,
           rowR_469,
           rowR_470,
           rowR_471,
           rowR_472,
           rowR_473,
           rowR_474,
           rowR_475,
           rowR_476,
           rowR_477,
           rowR_478,
           rowR_479,
           rowR_480,
           rowR_481,
           rowR_482,
           rowR_483,
           rowR_484,
           rowR_485,
           rowR_486,
           rowR_487,
           rowR_488,
           rowR_489,
           rowR_490,
           rowR_491,
           rowR_492,
           rowR_493,
           rowR_494,
           rowR_495,
           rowR_496,
           rowR_497,
           rowR_498,
           rowR_499,
           rowR_500,
           rowR_501,
           rowR_502,
           rowR_503,
           rowR_504,
           rowR_505,
           rowR_506,
           rowR_507,
           rowR_508,
           rowR_509,
           rowR_510,
           rowR_511,
           rowR_512,
           rowR_513,
           rowR_514,
           rowR_515,
           rowR_516,
           rowR_517,
           rowR_518,
           rowR_519,
           rowR_520,
           rowR_521,
           rowR_522,
           rowR_523,
           rowR_524,
           rowR_525,
           rowR_526,
           rowR_527,
           rowR_528,
           rowR_529,
           rowR_530,
           rowR_531,
           rowR_532,
           rowR_533,
           rowR_534,
           rowR_535,
           rowR_536,
           rowR_537,
           rowR_538,
           rowR_539,
           rowR_540,
           rowR_541,
           rowR_542,
           rowR_543,
           rowR_544,
           rowR_545,
           rowR_546,
           rowR_547,
           rowR_548,
           rowR_549,
           rowR_550,
           rowR_551,
           rowR_552,
           rowR_553,
           rowR_554,
           rowR_555,
           rowR_556,
           rowR_557,
           rowR_558,
           rowR_559,
           rowR_560,
           rowR_561,
           rowR_562,
           rowR_563,
           rowR_564,
           rowR_565,
           rowR_566,
           rowR_567,
           rowR_568,
           rowR_569,
           rowR_570,
           rowR_571,
           rowR_572,
           rowR_573,
           rowR_574,
           rowR_575,
           rowR_576,
           rowR_577,
           rowR_578,
           rowR_579,
           rowR_580,
           rowR_581,
           rowR_582,
           rowR_583,
           rowR_584,
           rowR_585,
           rowR_586,
           rowR_587,
           rowR_588,
           rowR_589,
           rowR_590,
           rowR_591,
           rowR_592,
           rowR_593,
           rowR_594,
           rowR_595,
           rowR_596,
           rowR_597,
           rowR_598,
           rowR_599,
           rowR_600,
           rowR_601,
           rowR_602,
           rowR_603,
           rowR_604,
           rowR_605,
           rowR_606,
           rowR_607,
           rowR_608,
           rowR_609,
           rowR_610,
           rowR_611,
           rowR_612,
           rowR_613,
           rowR_614,
           rowR_615,
           rowR_616,
           rowR_617,
           rowR_618,
           rowR_619,
           rowR_620,
           rowR_621,
           rowR_622,
           rowR_623,
           rowR_624,
           rowR_625,
           rowR_626,
           rowR_627,
           rowR_628,
           rowR_629,
           rowR_630,
           rowR_631,
           rowR_632,
           rowR_633,
           rowR_634,
           rowR_635,
           rowR_636,
           rowR_637,
           rowR_638,
           rowR_639,
           enS2P2
);

assign enC = enS2P1 & enS2P2;

Census_Transform_Row_fixpt census
          (clk,
          reset,
          clk_enable,
          rowL_0,
          rowL_1,
          rowL_2,
          rowL_3,
          rowL_4,
          rowL_5,
          rowL_6,
          rowL_7,
          rowL_8,
          rowL_9,
          rowL_10,
          rowL_11,
          rowL_12,
          rowL_13,
          rowL_14,
          rowL_15,
          rowL_16,
          rowL_17,
          rowL_18,
          rowL_19,
          rowL_20,
          rowL_21,
          rowL_22,
          rowL_23,
          rowL_24,
          rowL_25,
          rowL_26,
          rowL_27,
          rowL_28,
          rowL_29,
          rowL_30,
          rowL_31,
          rowL_32,
          rowL_33,
          rowL_34,
          rowL_35,
          rowL_36,
          rowL_37,
          rowL_38,
          rowL_39,
          rowL_40,
          rowL_41,
          rowL_42,
          rowL_43,
          rowL_44,
          rowL_45,
          rowL_46,
          rowL_47,
          rowL_48,
          rowL_49,
          rowL_50,
          rowL_51,
          rowL_52,
          rowL_53,
          rowL_54,
          rowL_55,
          rowL_56,
          rowL_57,
          rowL_58,
          rowL_59,
          rowL_60,
          rowL_61,
          rowL_62,
          rowL_63,
          rowL_64,
          rowL_65,
          rowL_66,
          rowL_67,
          rowL_68,
          rowL_69,
          rowL_70,
          rowL_71,
          rowL_72,
          rowL_73,
          rowL_74,
          rowL_75,
          rowL_76,
          rowL_77,
          rowL_78,
          rowL_79,
          rowL_80,
          rowL_81,
          rowL_82,
          rowL_83,
          rowL_84,
          rowL_85,
          rowL_86,
          rowL_87,
          rowL_88,
          rowL_89,
          rowL_90,
          rowL_91,
          rowL_92,
          rowL_93,
          rowL_94,
          rowL_95,
          rowL_96,
          rowL_97,
          rowL_98,
          rowL_99,
          rowL_100,
          rowL_101,
          rowL_102,
          rowL_103,
          rowL_104,
          rowL_105,
          rowL_106,
          rowL_107,
          rowL_108,
          rowL_109,
          rowL_110,
          rowL_111,
          rowL_112,
          rowL_113,
          rowL_114,
          rowL_115,
          rowL_116,
          rowL_117,
          rowL_118,
          rowL_119,
          rowL_120,
          rowL_121,
          rowL_122,
          rowL_123,
          rowL_124,
          rowL_125,
          rowL_126,
          rowL_127,
          rowL_128,
          rowL_129,
          rowL_130,
          rowL_131,
          rowL_132,
          rowL_133,
          rowL_134,
          rowL_135,
          rowL_136,
          rowL_137,
          rowL_138,
          rowL_139,
          rowL_140,
          rowL_141,
          rowL_142,
          rowL_143,
          rowL_144,
          rowL_145,
          rowL_146,
          rowL_147,
          rowL_148,
          rowL_149,
          rowL_150,
          rowL_151,
          rowL_152,
          rowL_153,
          rowL_154,
          rowL_155,
          rowL_156,
          rowL_157,
          rowL_158,
          rowL_159,
          rowL_160,
          rowL_161,
          rowL_162,
          rowL_163,
          rowL_164,
          rowL_165,
          rowL_166,
          rowL_167,
          rowL_168,
          rowL_169,
          rowL_170,
          rowL_171,
          rowL_172,
          rowL_173,
          rowL_174,
          rowL_175,
          rowL_176,
          rowL_177,
          rowL_178,
          rowL_179,
          rowL_180,
          rowL_181,
          rowL_182,
          rowL_183,
          rowL_184,
          rowL_185,
          rowL_186,
          rowL_187,
          rowL_188,
          rowL_189,
          rowL_190,
          rowL_191,
          rowL_192,
          rowL_193,
          rowL_194,
          rowL_195,
          rowL_196,
          rowL_197,
          rowL_198,
          rowL_199,
          rowL_200,
          rowL_201,
          rowL_202,
          rowL_203,
          rowL_204,
          rowL_205,
          rowL_206,
          rowL_207,
          rowL_208,
          rowL_209,
          rowL_210,
          rowL_211,
          rowL_212,
          rowL_213,
          rowL_214,
          rowL_215,
          rowL_216,
          rowL_217,
          rowL_218,
          rowL_219,
          rowL_220,
          rowL_221,
          rowL_222,
          rowL_223,
          rowL_224,
          rowL_225,
          rowL_226,
          rowL_227,
          rowL_228,
          rowL_229,
          rowL_230,
          rowL_231,
          rowL_232,
          rowL_233,
          rowL_234,
          rowL_235,
          rowL_236,
          rowL_237,
          rowL_238,
          rowL_239,
          rowL_240,
          rowL_241,
          rowL_242,
          rowL_243,
          rowL_244,
          rowL_245,
          rowL_246,
          rowL_247,
          rowL_248,
          rowL_249,
          rowL_250,
          rowL_251,
          rowL_252,
          rowL_253,
          rowL_254,
          rowL_255,
          rowL_256,
          rowL_257,
          rowL_258,
          rowL_259,
          rowL_260,
          rowL_261,
          rowL_262,
          rowL_263,
          rowL_264,
          rowL_265,
          rowL_266,
          rowL_267,
          rowL_268,
          rowL_269,
          rowL_270,
          rowL_271,
          rowL_272,
          rowL_273,
          rowL_274,
          rowL_275,
          rowL_276,
          rowL_277,
          rowL_278,
          rowL_279,
          rowL_280,
          rowL_281,
          rowL_282,
          rowL_283,
          rowL_284,
          rowL_285,
          rowL_286,
          rowL_287,
          rowL_288,
          rowL_289,
          rowL_290,
          rowL_291,
          rowL_292,
          rowL_293,
          rowL_294,
          rowL_295,
          rowL_296,
          rowL_297,
          rowL_298,
          rowL_299,
          rowL_300,
          rowL_301,
          rowL_302,
          rowL_303,
          rowL_304,
          rowL_305,
          rowL_306,
          rowL_307,
          rowL_308,
          rowL_309,
          rowL_310,
          rowL_311,
          rowL_312,
          rowL_313,
          rowL_314,
          rowL_315,
          rowL_316,
          rowL_317,
          rowL_318,
          rowL_319,
          rowL_320,
          rowL_321,
          rowL_322,
          rowL_323,
          rowL_324,
          rowL_325,
          rowL_326,
          rowL_327,
          rowL_328,
          rowL_329,
          rowL_330,
          rowL_331,
          rowL_332,
          rowL_333,
          rowL_334,
          rowL_335,
          rowL_336,
          rowL_337,
          rowL_338,
          rowL_339,
          rowL_340,
          rowL_341,
          rowL_342,
          rowL_343,
          rowL_344,
          rowL_345,
          rowL_346,
          rowL_347,
          rowL_348,
          rowL_349,
          rowL_350,
          rowL_351,
          rowL_352,
          rowL_353,
          rowL_354,
          rowL_355,
          rowL_356,
          rowL_357,
          rowL_358,
          rowL_359,
          rowL_360,
          rowL_361,
          rowL_362,
          rowL_363,
          rowL_364,
          rowL_365,
          rowL_366,
          rowL_367,
          rowL_368,
          rowL_369,
          rowL_370,
          rowL_371,
          rowL_372,
          rowL_373,
          rowL_374,
          rowL_375,
          rowL_376,
          rowL_377,
          rowL_378,
          rowL_379,
          rowL_380,
          rowL_381,
          rowL_382,
          rowL_383,
          rowL_384,
          rowL_385,
          rowL_386,
          rowL_387,
          rowL_388,
          rowL_389,
          rowL_390,
          rowL_391,
          rowL_392,
          rowL_393,
          rowL_394,
          rowL_395,
          rowL_396,
          rowL_397,
          rowL_398,
          rowL_399,
          rowL_400,
          rowL_401,
          rowL_402,
          rowL_403,
          rowL_404,
          rowL_405,
          rowL_406,
          rowL_407,
          rowL_408,
          rowL_409,
          rowL_410,
          rowL_411,
          rowL_412,
          rowL_413,
          rowL_414,
          rowL_415,
          rowL_416,
          rowL_417,
          rowL_418,
          rowL_419,
          rowL_420,
          rowL_421,
          rowL_422,
          rowL_423,
          rowL_424,
          rowL_425,
          rowL_426,
          rowL_427,
          rowL_428,
          rowL_429,
          rowL_430,
          rowL_431,
          rowL_432,
          rowL_433,
          rowL_434,
          rowL_435,
          rowL_436,
          rowL_437,
          rowL_438,
          rowL_439,
          rowL_440,
          rowL_441,
          rowL_442,
          rowL_443,
          rowL_444,
          rowL_445,
          rowL_446,
          rowL_447,
          rowL_448,
          rowL_449,
          rowL_450,
          rowL_451,
          rowL_452,
          rowL_453,
          rowL_454,
          rowL_455,
          rowL_456,
          rowL_457,
          rowL_458,
          rowL_459,
          rowL_460,
          rowL_461,
          rowL_462,
          rowL_463,
          rowL_464,
          rowL_465,
          rowL_466,
          rowL_467,
          rowL_468,
          rowL_469,
          rowL_470,
          rowL_471,
          rowL_472,
          rowL_473,
          rowL_474,
          rowL_475,
          rowL_476,
          rowL_477,
          rowL_478,
          rowL_479,
          rowL_480,
          rowL_481,
          rowL_482,
          rowL_483,
          rowL_484,
          rowL_485,
          rowL_486,
          rowL_487,
          rowL_488,
          rowL_489,
          rowL_490,
          rowL_491,
          rowL_492,
          rowL_493,
          rowL_494,
          rowL_495,
          rowL_496,
          rowL_497,
          rowL_498,
          rowL_499,
          rowL_500,
          rowL_501,
          rowL_502,
          rowL_503,
          rowL_504,
          rowL_505,
          rowL_506,
          rowL_507,
          rowL_508,
          rowL_509,
          rowL_510,
          rowL_511,
          rowL_512,
          rowL_513,
          rowL_514,
          rowL_515,
          rowL_516,
          rowL_517,
          rowL_518,
          rowL_519,
          rowL_520,
          rowL_521,
          rowL_522,
          rowL_523,
          rowL_524,
          rowL_525,
          rowL_526,
          rowL_527,
          rowL_528,
          rowL_529,
          rowL_530,
          rowL_531,
          rowL_532,
          rowL_533,
          rowL_534,
          rowL_535,
          rowL_536,
          rowL_537,
          rowL_538,
          rowL_539,
          rowL_540,
          rowL_541,
          rowL_542,
          rowL_543,
          rowL_544,
          rowL_545,
          rowL_546,
          rowL_547,
          rowL_548,
          rowL_549,
          rowL_550,
          rowL_551,
          rowL_552,
          rowL_553,
          rowL_554,
          rowL_555,
          rowL_556,
          rowL_557,
          rowL_558,
          rowL_559,
          rowL_560,
          rowL_561,
          rowL_562,
          rowL_563,
          rowL_564,
          rowL_565,
          rowL_566,
          rowL_567,
          rowL_568,
          rowL_569,
          rowL_570,
          rowL_571,
          rowL_572,
          rowL_573,
          rowL_574,
          rowL_575,
          rowL_576,
          rowL_577,
          rowL_578,
          rowL_579,
          rowL_580,
          rowL_581,
          rowL_582,
          rowL_583,
          rowL_584,
          rowL_585,
          rowL_586,
          rowL_587,
          rowL_588,
          rowL_589,
          rowL_590,
          rowL_591,
          rowL_592,
          rowL_593,
          rowL_594,
          rowL_595,
          rowL_596,
          rowL_597,
          rowL_598,
          rowL_599,
          rowL_600,
          rowL_601,
          rowL_602,
          rowL_603,
          rowL_604,
          rowL_605,
          rowL_606,
          rowL_607,
          rowL_608,
          rowL_609,
          rowL_610,
          rowL_611,
          rowL_612,
          rowL_613,
          rowL_614,
          rowL_615,
          rowL_616,
          rowL_617,
          rowL_618,
          rowL_619,
          rowL_620,
          rowL_621,
          rowL_622,
          rowL_623,
          rowL_624,
          rowL_625,
          rowL_626,
          rowL_627,
          rowL_628,
          rowL_629,
          rowL_630,
          rowL_631,
          rowL_632,
          rowL_633,
          rowL_634,
          rowL_635,
          rowL_636,
          rowL_637,
          rowL_638,
          rowL_639,           
          rowR_0,
          rowR_1,
          rowR_2,
          rowR_3,
          rowR_4,
          rowR_5,
          rowR_6,
          rowR_7,
          rowR_8,
          rowR_9,
          rowR_10,
          rowR_11,
          rowR_12,
          rowR_13,
          rowR_14,
          rowR_15,
          rowR_16,
          rowR_17,
          rowR_18,
          rowR_19,
          rowR_20,
          rowR_21,
          rowR_22,
          rowR_23,
          rowR_24,
          rowR_25,
          rowR_26,
          rowR_27,
          rowR_28,
          rowR_29,
          rowR_30,
          rowR_31,
          rowR_32,
          rowR_33,
          rowR_34,
          rowR_35,
          rowR_36,
          rowR_37,
          rowR_38,
          rowR_39,
          rowR_40,
          rowR_41,
          rowR_42,
          rowR_43,
          rowR_44,
          rowR_45,
          rowR_46,
          rowR_47,
          rowR_48,
          rowR_49,
          rowR_50,
          rowR_51,
          rowR_52,
          rowR_53,
          rowR_54,
          rowR_55,
          rowR_56,
          rowR_57,
          rowR_58,
          rowR_59,
          rowR_60,
          rowR_61,
          rowR_62,
          rowR_63,
          rowR_64,
          rowR_65,
          rowR_66,
          rowR_67,
          rowR_68,
          rowR_69,
          rowR_70,
          rowR_71,
          rowR_72,
          rowR_73,
          rowR_74,
          rowR_75,
          rowR_76,
          rowR_77,
          rowR_78,
          rowR_79,
          rowR_80,
          rowR_81,
          rowR_82,
          rowR_83,
          rowR_84,
          rowR_85,
          rowR_86,
          rowR_87,
          rowR_88,
          rowR_89,
          rowR_90,
          rowR_91,
          rowR_92,
          rowR_93,
          rowR_94,
          rowR_95,
          rowR_96,
          rowR_97,
          rowR_98,
          rowR_99,
          rowR_100,
          rowR_101,
          rowR_102,
          rowR_103,
          rowR_104,
          rowR_105,
          rowR_106,
          rowR_107,
          rowR_108,
          rowR_109,
          rowR_110,
          rowR_111,
          rowR_112,
          rowR_113,
          rowR_114,
          rowR_115,
          rowR_116,
          rowR_117,
          rowR_118,
          rowR_119,
          rowR_120,
          rowR_121,
          rowR_122,
          rowR_123,
          rowR_124,
          rowR_125,
          rowR_126,
          rowR_127,
          rowR_128,
          rowR_129,
          rowR_130,
          rowR_131,
          rowR_132,
          rowR_133,
          rowR_134,
          rowR_135,
          rowR_136,
          rowR_137,
          rowR_138,
          rowR_139,
          rowR_140,
          rowR_141,
          rowR_142,
          rowR_143,
          rowR_144,
          rowR_145,
          rowR_146,
          rowR_147,
          rowR_148,
          rowR_149,
          rowR_150,
          rowR_151,
          rowR_152,
          rowR_153,
          rowR_154,
          rowR_155,
          rowR_156,
          rowR_157,
          rowR_158,
          rowR_159,
          rowR_160,
          rowR_161,
          rowR_162,
          rowR_163,
          rowR_164,
          rowR_165,
          rowR_166,
          rowR_167,
          rowR_168,
          rowR_169,
          rowR_170,
          rowR_171,
          rowR_172,
          rowR_173,
          rowR_174,
          rowR_175,
          rowR_176,
          rowR_177,
          rowR_178,
          rowR_179,
          rowR_180,
          rowR_181,
          rowR_182,
          rowR_183,
          rowR_184,
          rowR_185,
          rowR_186,
          rowR_187,
          rowR_188,
          rowR_189,
          rowR_190,
          rowR_191,
          rowR_192,
          rowR_193,
          rowR_194,
          rowR_195,
          rowR_196,
          rowR_197,
          rowR_198,
          rowR_199,
          rowR_200,
          rowR_201,
          rowR_202,
          rowR_203,
          rowR_204,
          rowR_205,
          rowR_206,
          rowR_207,
          rowR_208,
          rowR_209,
          rowR_210,
          rowR_211,
          rowR_212,
          rowR_213,
          rowR_214,
          rowR_215,
          rowR_216,
          rowR_217,
          rowR_218,
          rowR_219,
          rowR_220,
          rowR_221,
          rowR_222,
          rowR_223,
          rowR_224,
          rowR_225,
          rowR_226,
          rowR_227,
          rowR_228,
          rowR_229,
          rowR_230,
          rowR_231,
          rowR_232,
          rowR_233,
          rowR_234,
          rowR_235,
          rowR_236,
          rowR_237,
          rowR_238,
          rowR_239,
          rowR_240,
          rowR_241,
          rowR_242,
          rowR_243,
          rowR_244,
          rowR_245,
          rowR_246,
          rowR_247,
          rowR_248,
          rowR_249,
          rowR_250,
          rowR_251,
          rowR_252,
          rowR_253,
          rowR_254,
          rowR_255,
          rowR_256,
          rowR_257,
          rowR_258,
          rowR_259,
          rowR_260,
          rowR_261,
          rowR_262,
          rowR_263,
          rowR_264,
          rowR_265,
          rowR_266,
          rowR_267,
          rowR_268,
          rowR_269,
          rowR_270,
          rowR_271,
          rowR_272,
          rowR_273,
          rowR_274,
          rowR_275,
          rowR_276,
          rowR_277,
          rowR_278,
          rowR_279,
          rowR_280,
          rowR_281,
          rowR_282,
          rowR_283,
          rowR_284,
          rowR_285,
          rowR_286,
          rowR_287,
          rowR_288,
          rowR_289,
          rowR_290,
          rowR_291,
          rowR_292,
          rowR_293,
          rowR_294,
          rowR_295,
          rowR_296,
          rowR_297,
          rowR_298,
          rowR_299,
          rowR_300,
          rowR_301,
          rowR_302,
          rowR_303,
          rowR_304,
          rowR_305,
          rowR_306,
          rowR_307,
          rowR_308,
          rowR_309,
          rowR_310,
          rowR_311,
          rowR_312,
          rowR_313,
          rowR_314,
          rowR_315,
          rowR_316,
          rowR_317,
          rowR_318,
          rowR_319,
          rowR_320,
          rowR_321,
          rowR_322,
          rowR_323,
          rowR_324,
          rowR_325,
          rowR_326,
          rowR_327,
          rowR_328,
          rowR_329,
          rowR_330,
          rowR_331,
          rowR_332,
          rowR_333,
          rowR_334,
          rowR_335,
          rowR_336,
          rowR_337,
          rowR_338,
          rowR_339,
          rowR_340,
          rowR_341,
          rowR_342,
          rowR_343,
          rowR_344,
          rowR_345,
          rowR_346,
          rowR_347,
          rowR_348,
          rowR_349,
          rowR_350,
          rowR_351,
          rowR_352,
          rowR_353,
          rowR_354,
          rowR_355,
          rowR_356,
          rowR_357,
          rowR_358,
          rowR_359,
          rowR_360,
          rowR_361,
          rowR_362,
          rowR_363,
          rowR_364,
          rowR_365,
          rowR_366,
          rowR_367,
          rowR_368,
          rowR_369,
          rowR_370,
          rowR_371,
          rowR_372,
          rowR_373,
          rowR_374,
          rowR_375,
          rowR_376,
          rowR_377,
          rowR_378,
          rowR_379,
          rowR_380,
          rowR_381,
          rowR_382,
          rowR_383,
          rowR_384,
          rowR_385,
          rowR_386,
          rowR_387,
          rowR_388,
          rowR_389,
          rowR_390,
          rowR_391,
          rowR_392,
          rowR_393,
          rowR_394,
          rowR_395,
          rowR_396,
          rowR_397,
          rowR_398,
          rowR_399,
          rowR_400,
          rowR_401,
          rowR_402,
          rowR_403,
          rowR_404,
          rowR_405,
          rowR_406,
          rowR_407,
          rowR_408,
          rowR_409,
          rowR_410,
          rowR_411,
          rowR_412,
          rowR_413,
          rowR_414,
          rowR_415,
          rowR_416,
          rowR_417,
          rowR_418,
          rowR_419,
          rowR_420,
          rowR_421,
          rowR_422,
          rowR_423,
          rowR_424,
          rowR_425,
          rowR_426,
          rowR_427,
          rowR_428,
          rowR_429,
          rowR_430,
          rowR_431,
          rowR_432,
          rowR_433,
          rowR_434,
          rowR_435,
          rowR_436,
          rowR_437,
          rowR_438,
          rowR_439,
          rowR_440,
          rowR_441,
          rowR_442,
          rowR_443,
          rowR_444,
          rowR_445,
          rowR_446,
          rowR_447,
          rowR_448,
          rowR_449,
          rowR_450,
          rowR_451,
          rowR_452,
          rowR_453,
          rowR_454,
          rowR_455,
          rowR_456,
          rowR_457,
          rowR_458,
          rowR_459,
          rowR_460,
          rowR_461,
          rowR_462,
          rowR_463,
          rowR_464,
          rowR_465,
          rowR_466,
          rowR_467,
          rowR_468,
          rowR_469,
          rowR_470,
          rowR_471,
          rowR_472,
          rowR_473,
          rowR_474,
          rowR_475,
          rowR_476,
          rowR_477,
          rowR_478,
          rowR_479,
          rowR_480,
          rowR_481,
          rowR_482,
          rowR_483,
          rowR_484,
          rowR_485,
          rowR_486,
          rowR_487,
          rowR_488,
          rowR_489,
          rowR_490,
          rowR_491,
          rowR_492,
          rowR_493,
          rowR_494,
          rowR_495,
          rowR_496,
          rowR_497,
          rowR_498,
          rowR_499,
          rowR_500,
          rowR_501,
          rowR_502,
          rowR_503,
          rowR_504,
          rowR_505,
          rowR_506,
          rowR_507,
          rowR_508,
          rowR_509,
          rowR_510,
          rowR_511,
          rowR_512,
          rowR_513,
          rowR_514,
          rowR_515,
          rowR_516,
          rowR_517,
          rowR_518,
          rowR_519,
          rowR_520,
          rowR_521,
          rowR_522,
          rowR_523,
          rowR_524,
          rowR_525,
          rowR_526,
          rowR_527,
          rowR_528,
          rowR_529,
          rowR_530,
          rowR_531,
          rowR_532,
          rowR_533,
          rowR_534,
          rowR_535,
          rowR_536,
          rowR_537,
          rowR_538,
          rowR_539,
          rowR_540,
          rowR_541,
          rowR_542,
          rowR_543,
          rowR_544,
          rowR_545,
          rowR_546,
          rowR_547,
          rowR_548,
          rowR_549,
          rowR_550,
          rowR_551,
          rowR_552,
          rowR_553,
          rowR_554,
          rowR_555,
          rowR_556,
          rowR_557,
          rowR_558,
          rowR_559,
          rowR_560,
          rowR_561,
          rowR_562,
          rowR_563,
          rowR_564,
          rowR_565,
          rowR_566,
          rowR_567,
          rowR_568,
          rowR_569,
          rowR_570,
          rowR_571,
          rowR_572,
          rowR_573,
          rowR_574,
          rowR_575,
          rowR_576,
          rowR_577,
          rowR_578,
          rowR_579,
          rowR_580,
          rowR_581,
          rowR_582,
          rowR_583,
          rowR_584,
          rowR_585,
          rowR_586,
          rowR_587,
          rowR_588,
          rowR_589,
          rowR_590,
          rowR_591,
          rowR_592,
          rowR_593,
          rowR_594,
          rowR_595,
          rowR_596,
          rowR_597,
          rowR_598,
          rowR_599,
          rowR_600,
          rowR_601,
          rowR_602,
          rowR_603,
          rowR_604,
          rowR_605,
          rowR_606,
          rowR_607,
          rowR_608,
          rowR_609,
          rowR_610,
          rowR_611,
          rowR_612,
          rowR_613,
          rowR_614,
          rowR_615,
          rowR_616,
          rowR_617,
          rowR_618,
          rowR_619,
          rowR_620,
          rowR_621,
          rowR_622,
          rowR_623,
          rowR_624,
          rowR_625,
          rowR_626,
          rowR_627,
          rowR_628,
          rowR_629,
          rowR_630,
          rowR_631,
          rowR_632,
          rowR_633,
          rowR_634,
          rowR_635,
          rowR_636,
          rowR_637,
          rowR_638,
          rowR_639,
          enC,
          ce_out3,
          rowD_0,
          rowD_1,
          rowD_2,
          rowD_3,
          rowD_4,
          rowD_5,
          rowD_6,
          rowD_7,
          rowD_8,
          rowD_9,
          rowD_10,
          rowD_11,
          rowD_12,
          rowD_13,
          rowD_14,
          rowD_15,
          rowD_16,
          rowD_17,
          rowD_18,
          rowD_19,
          rowD_20,
          rowD_21,
          rowD_22,
          rowD_23,
          rowD_24,
          rowD_25,
          rowD_26,
          rowD_27,
          rowD_28,
          rowD_29,
          rowD_30,
          rowD_31,
          rowD_32,
          rowD_33,
          rowD_34,
          rowD_35,
          rowD_36,
          rowD_37,
          rowD_38,
          rowD_39,
          rowD_40,
          rowD_41,
          rowD_42,
          rowD_43,
          rowD_44,
          rowD_45,
          rowD_46,
          rowD_47,
          rowD_48,
          rowD_49,
          rowD_50,
          rowD_51,
          rowD_52,
          rowD_53,
          rowD_54,
          rowD_55,
          rowD_56,
          rowD_57,
          rowD_58,
          rowD_59,
          rowD_60,
          rowD_61,
          rowD_62,
          rowD_63,
          rowD_64,
          rowD_65,
          rowD_66,
          rowD_67,
          rowD_68,
          rowD_69,
          rowD_70,
          rowD_71,
          rowD_72,
          rowD_73,
          rowD_74,
          rowD_75,
          rowD_76,
          rowD_77,
          rowD_78,
          rowD_79,
          rowD_80,
          rowD_81,
          rowD_82,
          rowD_83,
          rowD_84,
          rowD_85,
          rowD_86,
          rowD_87,
          rowD_88,
          rowD_89,
          rowD_90,
          rowD_91,
          rowD_92,
          rowD_93,
          rowD_94,
          rowD_95,
          rowD_96,
          rowD_97,
          rowD_98,
          rowD_99,
          rowD_100,
          rowD_101,
          rowD_102,
          rowD_103,
          rowD_104,
          rowD_105,
          rowD_106,
          rowD_107,
          rowD_108,
          rowD_109,
          rowD_110,
          rowD_111,
          rowD_112,
          rowD_113,
          rowD_114,
          rowD_115,
          rowD_116,
          rowD_117,
          rowD_118,
          rowD_119,
          rowD_120,
          rowD_121,
          rowD_122,
          rowD_123,
          rowD_124,
          rowD_125,
          rowD_126,
          rowD_127,
          rowD_128,
          rowD_129,
          rowD_130,
          rowD_131,
          rowD_132,
          rowD_133,
          rowD_134,
          rowD_135,
          rowD_136,
          rowD_137,
          rowD_138,
          rowD_139,
          rowD_140,
          rowD_141,
          rowD_142,
          rowD_143,
          rowD_144,
          rowD_145,
          rowD_146,
          rowD_147,
          rowD_148,
          rowD_149,
          rowD_150,
          rowD_151,
          rowD_152,
          rowD_153,
          rowD_154,
          rowD_155,
          rowD_156,
          rowD_157,
          rowD_158,
          rowD_159,
          rowD_160,
          rowD_161,
          rowD_162,
          rowD_163,
          rowD_164,
          rowD_165,
          rowD_166,
          rowD_167,
          rowD_168,
          rowD_169,
          rowD_170,
          rowD_171,
          rowD_172,
          rowD_173,
          rowD_174,
          rowD_175,
          rowD_176,
          rowD_177,
          rowD_178,
          rowD_179,
          rowD_180,
          rowD_181,
          rowD_182,
          rowD_183,
          rowD_184,
          rowD_185,
          rowD_186,
          rowD_187,
          rowD_188,
          rowD_189,
          rowD_190,
          rowD_191,
          rowD_192,
          rowD_193,
          rowD_194,
          rowD_195,
          rowD_196,
          rowD_197,
          rowD_198,
          rowD_199,
          rowD_200,
          rowD_201,
          rowD_202,
          rowD_203,
          rowD_204,
          rowD_205,
          rowD_206,
          rowD_207,
          rowD_208,
          rowD_209,
          rowD_210,
          rowD_211,
          rowD_212,
          rowD_213,
          rowD_214,
          rowD_215,
          rowD_216,
          rowD_217,
          rowD_218,
          rowD_219,
          rowD_220,
          rowD_221,
          rowD_222,
          rowD_223,
          rowD_224,
          rowD_225,
          rowD_226,
          rowD_227,
          rowD_228,
          rowD_229,
          rowD_230,
          rowD_231,
          rowD_232,
          rowD_233,
          rowD_234,
          rowD_235,
          rowD_236,
          rowD_237,
          rowD_238,
          rowD_239,
          rowD_240,
          rowD_241,
          rowD_242,
          rowD_243,
          rowD_244,
          rowD_245,
          rowD_246,
          rowD_247,
          rowD_248,
          rowD_249,
          rowD_250,
          rowD_251,
          rowD_252,
          rowD_253,
          rowD_254,
          rowD_255,
          rowD_256,
          rowD_257,
          rowD_258,
          rowD_259,
          rowD_260,
          rowD_261,
          rowD_262,
          rowD_263,
          rowD_264,
          rowD_265,
          rowD_266,
          rowD_267,
          rowD_268,
          rowD_269,
          rowD_270,
          rowD_271,
          rowD_272,
          rowD_273,
          rowD_274,
          rowD_275,
          rowD_276,
          rowD_277,
          rowD_278,
          rowD_279,
          rowD_280,
          rowD_281,
          rowD_282,
          rowD_283,
          rowD_284,
          rowD_285,
          rowD_286,
          rowD_287,
          rowD_288,
          rowD_289,
          rowD_290,
          rowD_291,
          rowD_292,
          rowD_293,
          rowD_294,
          rowD_295,
          rowD_296,
          rowD_297,
          rowD_298,
          rowD_299,
          rowD_300,
          rowD_301,
          rowD_302,
          rowD_303,
          rowD_304,
          rowD_305,
          rowD_306,
          rowD_307,
          rowD_308,
          rowD_309,
          rowD_310,
          rowD_311,
          rowD_312,
          rowD_313,
          rowD_314,
          rowD_315,
          rowD_316,
          rowD_317,
          rowD_318,
          rowD_319,
          rowD_320,
          rowD_321,
          rowD_322,
          rowD_323,
          rowD_324,
          rowD_325,
          rowD_326,
          rowD_327,
          rowD_328,
          rowD_329,
          rowD_330,
          rowD_331,
          rowD_332,
          rowD_333,
          rowD_334,
          rowD_335,
          rowD_336,
          rowD_337,
          rowD_338,
          rowD_339,
          rowD_340,
          rowD_341,
          rowD_342,
          rowD_343,
          rowD_344,
          rowD_345,
          rowD_346,
          rowD_347,
          rowD_348,
          rowD_349,
          rowD_350,
          rowD_351,
          rowD_352,
          rowD_353,
          rowD_354,
          rowD_355,
          rowD_356,
          rowD_357,
          rowD_358,
          rowD_359,
          rowD_360,
          rowD_361,
          rowD_362,
          rowD_363,
          rowD_364,
          rowD_365,
          rowD_366,
          rowD_367,
          rowD_368,
          rowD_369,
          rowD_370,
          rowD_371,
          rowD_372,
          rowD_373,
          rowD_374,
          rowD_375,
          rowD_376,
          rowD_377,
          rowD_378,
          rowD_379,
          rowD_380,
          rowD_381,
          rowD_382,
          rowD_383,
          rowD_384,
          rowD_385,
          rowD_386,
          rowD_387,
          rowD_388,
          rowD_389,
          rowD_390,
          rowD_391,
          rowD_392,
          rowD_393,
          rowD_394,
          rowD_395,
          rowD_396,
          rowD_397,
          rowD_398,
          rowD_399,
          rowD_400,
          rowD_401,
          rowD_402,
          rowD_403,
          rowD_404,
          rowD_405,
          rowD_406,
          rowD_407,
          rowD_408,
          rowD_409,
          rowD_410,
          rowD_411,
          rowD_412,
          rowD_413,
          rowD_414,
          rowD_415,
          rowD_416,
          rowD_417,
          rowD_418,
          rowD_419,
          rowD_420,
          rowD_421,
          rowD_422,
          rowD_423,
          rowD_424,
          rowD_425,
          rowD_426,
          rowD_427,
          rowD_428,
          rowD_429,
          rowD_430,
          rowD_431,
          rowD_432,
          rowD_433,
          rowD_434,
          rowD_435,
          rowD_436,
          rowD_437,
          rowD_438,
          rowD_439,
          rowD_440,
          rowD_441,
          rowD_442,
          rowD_443,
          rowD_444,
          rowD_445,
          rowD_446,
          rowD_447,
          rowD_448,
          rowD_449,
          rowD_450,
          rowD_451,
          rowD_452,
          rowD_453,
          rowD_454,
          rowD_455,
          rowD_456,
          rowD_457,
          rowD_458,
          rowD_459,
          rowD_460,
          rowD_461,
          rowD_462,
          rowD_463,
          rowD_464,
          rowD_465,
          rowD_466,
          rowD_467,
          rowD_468,
          rowD_469,
          rowD_470,
          rowD_471,
          rowD_472,
          rowD_473,
          rowD_474,
          rowD_475,
          rowD_476,
          rowD_477,
          rowD_478,
          rowD_479,
          rowD_480,
          rowD_481,
          rowD_482,
          rowD_483,
          rowD_484,
          rowD_485,
          rowD_486,
          rowD_487,
          rowD_488,
          rowD_489,
          rowD_490,
          rowD_491,
          rowD_492,
          rowD_493,
          rowD_494,
          rowD_495,
          rowD_496,
          rowD_497,
          rowD_498,
          rowD_499,
          rowD_500,
          rowD_501,
          rowD_502,
          rowD_503,
          rowD_504,
          rowD_505,
          rowD_506,
          rowD_507,
          rowD_508,
          rowD_509,
          rowD_510,
          rowD_511,
          rowD_512,
          rowD_513,
          rowD_514,
          rowD_515,
          rowD_516,
          rowD_517,
          rowD_518,
          rowD_519,
          rowD_520,
          rowD_521,
          rowD_522,
          rowD_523,
          rowD_524,
          rowD_525,
          rowD_526,
          rowD_527,
          rowD_528,
          rowD_529,
          rowD_530,
          rowD_531,
          rowD_532,
          rowD_533,
          rowD_534,
          rowD_535,
          rowD_536,
          rowD_537,
          rowD_538,
          rowD_539,
          rowD_540,
          rowD_541,
          rowD_542,
          rowD_543,
          rowD_544,
          rowD_545,
          rowD_546,
          rowD_547,
          rowD_548,
          rowD_549,
          rowD_550,
          rowD_551,
          rowD_552,
          rowD_553,
          rowD_554,
          rowD_555,
          rowD_556,
          rowD_557,
          rowD_558,
          rowD_559,
          rowD_560,
          rowD_561,
          rowD_562,
          rowD_563,
          rowD_564,
          rowD_565,
          rowD_566,
          rowD_567,
          rowD_568,
          rowD_569,
          rowD_570,
          rowD_571,
          rowD_572,
          rowD_573,
          rowD_574,
          rowD_575,
          rowD_576,
          rowD_577,
          rowD_578,
          rowD_579,
          rowD_580,
          rowD_581,
          rowD_582,
          rowD_583,
          rowD_584,
          rowD_585,
          rowD_586,
          rowD_587,
          rowD_588,
          rowD_589,
          rowD_590,
          rowD_591,
          rowD_592,
          rowD_593,
          rowD_594,
          rowD_595,
          rowD_596,
          rowD_597,
          rowD_598,
          rowD_599,
          rowD_600,
          rowD_601,
          rowD_602,
          rowD_603,
          rowD_604,
          rowD_605,
          rowD_606,
          rowD_607,
          rowD_608,
          rowD_609,
          rowD_610,
          rowD_611,
          rowD_612,
          rowD_613,
          rowD_614,
          rowD_615,
          rowD_616,
          rowD_617,
          rowD_618,
          rowD_619,
          rowD_620,
          rowD_621,
          rowD_622,
          rowD_623,
          rowD_624,
          rowD_625,
          rowD_626,
          rowD_627,
          rowD_628,
          rowD_629,
          rowD_630,
          rowD_631,
          rowD_632,
          rowD_633,
          rowD_634,
          rowD_635,
          rowD_636,
          rowD_637,
          rowD_638,
          rowD_639,
          enP2S
);

Parallel_to_Serial_fixpt ps1
         (clk,
         reset,
         clk_enable,
         rowD_0,
         rowD_1,
         rowD_2,
         rowD_3,
         rowD_4,
         rowD_5,
         rowD_6,
         rowD_7,
         rowD_8,
         rowD_9,
         rowD_10,
         rowD_11,
         rowD_12,
         rowD_13,
         rowD_14,
         rowD_15,
         rowD_16,
         rowD_17,
         rowD_18,
         rowD_19,
         rowD_20,
         rowD_21,
         rowD_22,
         rowD_23,
         rowD_24,
         rowD_25,
         rowD_26,
         rowD_27,
         rowD_28,
         rowD_29,
         rowD_30,
         rowD_31,
         rowD_32,
         rowD_33,
         rowD_34,
         rowD_35,
         rowD_36,
         rowD_37,
         rowD_38,
         rowD_39,
         rowD_40,
         rowD_41,
         rowD_42,
         rowD_43,
         rowD_44,
         rowD_45,
         rowD_46,
         rowD_47,
         rowD_48,
         rowD_49,
         rowD_50,
         rowD_51,
         rowD_52,
         rowD_53,
         rowD_54,
         rowD_55,
         rowD_56,
         rowD_57,
         rowD_58,
         rowD_59,
         rowD_60,
         rowD_61,
         rowD_62,
         rowD_63,
         rowD_64,
         rowD_65,
         rowD_66,
         rowD_67,
         rowD_68,
         rowD_69,
         rowD_70,
         rowD_71,
         rowD_72,
         rowD_73,
         rowD_74,
         rowD_75,
         rowD_76,
         rowD_77,
         rowD_78,
         rowD_79,
         rowD_80,
         rowD_81,
         rowD_82,
         rowD_83,
         rowD_84,
         rowD_85,
         rowD_86,
         rowD_87,
         rowD_88,
         rowD_89,
         rowD_90,
         rowD_91,
         rowD_92,
         rowD_93,
         rowD_94,
         rowD_95,
         rowD_96,
         rowD_97,
         rowD_98,
         rowD_99,
         rowD_100,
         rowD_101,
         rowD_102,
         rowD_103,
         rowD_104,
         rowD_105,
         rowD_106,
         rowD_107,
         rowD_108,
         rowD_109,
         rowD_110,
         rowD_111,
         rowD_112,
         rowD_113,
         rowD_114,
         rowD_115,
         rowD_116,
         rowD_117,
         rowD_118,
         rowD_119,
         rowD_120,
         rowD_121,
         rowD_122,
         rowD_123,
         rowD_124,
         rowD_125,
         rowD_126,
         rowD_127,
         rowD_128,
         rowD_129,
         rowD_130,
         rowD_131,
         rowD_132,
         rowD_133,
         rowD_134,
         rowD_135,
         rowD_136,
         rowD_137,
         rowD_138,
         rowD_139,
         rowD_140,
         rowD_141,
         rowD_142,
         rowD_143,
         rowD_144,
         rowD_145,
         rowD_146,
         rowD_147,
         rowD_148,
         rowD_149,
         rowD_150,
         rowD_151,
         rowD_152,
         rowD_153,
         rowD_154,
         rowD_155,
         rowD_156,
         rowD_157,
         rowD_158,
         rowD_159,
         rowD_160,
         rowD_161,
         rowD_162,
         rowD_163,
         rowD_164,
         rowD_165,
         rowD_166,
         rowD_167,
         rowD_168,
         rowD_169,
         rowD_170,
         rowD_171,
         rowD_172,
         rowD_173,
         rowD_174,
         rowD_175,
         rowD_176,
         rowD_177,
         rowD_178,
         rowD_179,
         rowD_180,
         rowD_181,
         rowD_182,
         rowD_183,
         rowD_184,
         rowD_185,
         rowD_186,
         rowD_187,
         rowD_188,
         rowD_189,
         rowD_190,
         rowD_191,
         rowD_192,
         rowD_193,
         rowD_194,
         rowD_195,
         rowD_196,
         rowD_197,
         rowD_198,
         rowD_199,
         rowD_200,
         rowD_201,
         rowD_202,
         rowD_203,
         rowD_204,
         rowD_205,
         rowD_206,
         rowD_207,
         rowD_208,
         rowD_209,
         rowD_210,
         rowD_211,
         rowD_212,
         rowD_213,
         rowD_214,
         rowD_215,
         rowD_216,
         rowD_217,
         rowD_218,
         rowD_219,
         rowD_220,
         rowD_221,
         rowD_222,
         rowD_223,
         rowD_224,
         rowD_225,
         rowD_226,
         rowD_227,
         rowD_228,
         rowD_229,
         rowD_230,
         rowD_231,
         rowD_232,
         rowD_233,
         rowD_234,
         rowD_235,
         rowD_236,
         rowD_237,
         rowD_238,
         rowD_239,
         rowD_240,
         rowD_241,
         rowD_242,
         rowD_243,
         rowD_244,
         rowD_245,
         rowD_246,
         rowD_247,
         rowD_248,
         rowD_249,
         rowD_250,
         rowD_251,
         rowD_252,
         rowD_253,
         rowD_254,
         rowD_255,
         rowD_256,
         rowD_257,
         rowD_258,
         rowD_259,
         rowD_260,
         rowD_261,
         rowD_262,
         rowD_263,
         rowD_264,
         rowD_265,
         rowD_266,
         rowD_267,
         rowD_268,
         rowD_269,
         rowD_270,
         rowD_271,
         rowD_272,
         rowD_273,
         rowD_274,
         rowD_275,
         rowD_276,
         rowD_277,
         rowD_278,
         rowD_279,
         rowD_280,
         rowD_281,
         rowD_282,
         rowD_283,
         rowD_284,
         rowD_285,
         rowD_286,
         rowD_287,
         rowD_288,
         rowD_289,
         rowD_290,
         rowD_291,
         rowD_292,
         rowD_293,
         rowD_294,
         rowD_295,
         rowD_296,
         rowD_297,
         rowD_298,
         rowD_299,
         rowD_300,
         rowD_301,
         rowD_302,
         rowD_303,
         rowD_304,
         rowD_305,
         rowD_306,
         rowD_307,
         rowD_308,
         rowD_309,
         rowD_310,
         rowD_311,
         rowD_312,
         rowD_313,
         rowD_314,
         rowD_315,
         rowD_316,
         rowD_317,
         rowD_318,
         rowD_319,
         rowD_320,
         rowD_321,
         rowD_322,
         rowD_323,
         rowD_324,
         rowD_325,
         rowD_326,
         rowD_327,
         rowD_328,
         rowD_329,
         rowD_330,
         rowD_331,
         rowD_332,
         rowD_333,
         rowD_334,
         rowD_335,
         rowD_336,
         rowD_337,
         rowD_338,
         rowD_339,
         rowD_340,
         rowD_341,
         rowD_342,
         rowD_343,
         rowD_344,
         rowD_345,
         rowD_346,
         rowD_347,
         rowD_348,
         rowD_349,
         rowD_350,
         rowD_351,
         rowD_352,
         rowD_353,
         rowD_354,
         rowD_355,
         rowD_356,
         rowD_357,
         rowD_358,
         rowD_359,
         rowD_360,
         rowD_361,
         rowD_362,
         rowD_363,
         rowD_364,
         rowD_365,
         rowD_366,
         rowD_367,
         rowD_368,
         rowD_369,
         rowD_370,
         rowD_371,
         rowD_372,
         rowD_373,
         rowD_374,
         rowD_375,
         rowD_376,
         rowD_377,
         rowD_378,
         rowD_379,
         rowD_380,
         rowD_381,
         rowD_382,
         rowD_383,
         rowD_384,
         rowD_385,
         rowD_386,
         rowD_387,
         rowD_388,
         rowD_389,
         rowD_390,
         rowD_391,
         rowD_392,
         rowD_393,
         rowD_394,
         rowD_395,
         rowD_396,
         rowD_397,
         rowD_398,
         rowD_399,
         rowD_400,
         rowD_401,
         rowD_402,
         rowD_403,
         rowD_404,
         rowD_405,
         rowD_406,
         rowD_407,
         rowD_408,
         rowD_409,
         rowD_410,
         rowD_411,
         rowD_412,
         rowD_413,
         rowD_414,
         rowD_415,
         rowD_416,
         rowD_417,
         rowD_418,
         rowD_419,
         rowD_420,
         rowD_421,
         rowD_422,
         rowD_423,
         rowD_424,
         rowD_425,
         rowD_426,
         rowD_427,
         rowD_428,
         rowD_429,
         rowD_430,
         rowD_431,
         rowD_432,
         rowD_433,
         rowD_434,
         rowD_435,
         rowD_436,
         rowD_437,
         rowD_438,
         rowD_439,
         rowD_440,
         rowD_441,
         rowD_442,
         rowD_443,
         rowD_444,
         rowD_445,
         rowD_446,
         rowD_447,
         rowD_448,
         rowD_449,
         rowD_450,
         rowD_451,
         rowD_452,
         rowD_453,
         rowD_454,
         rowD_455,
         rowD_456,
         rowD_457,
         rowD_458,
         rowD_459,
         rowD_460,
         rowD_461,
         rowD_462,
         rowD_463,
         rowD_464,
         rowD_465,
         rowD_466,
         rowD_467,
         rowD_468,
         rowD_469,
         rowD_470,
         rowD_471,
         rowD_472,
         rowD_473,
         rowD_474,
         rowD_475,
         rowD_476,
         rowD_477,
         rowD_478,
         rowD_479,
         rowD_480,
         rowD_481,
         rowD_482,
         rowD_483,
         rowD_484,
         rowD_485,
         rowD_486,
         rowD_487,
         rowD_488,
         rowD_489,
         rowD_490,
         rowD_491,
         rowD_492,
         rowD_493,
         rowD_494,
         rowD_495,
         rowD_496,
         rowD_497,
         rowD_498,
         rowD_499,
         rowD_500,
         rowD_501,
         rowD_502,
         rowD_503,
         rowD_504,
         rowD_505,
         rowD_506,
         rowD_507,
         rowD_508,
         rowD_509,
         rowD_510,
         rowD_511,
         rowD_512,
         rowD_513,
         rowD_514,
         rowD_515,
         rowD_516,
         rowD_517,
         rowD_518,
         rowD_519,
         rowD_520,
         rowD_521,
         rowD_522,
         rowD_523,
         rowD_524,
         rowD_525,
         rowD_526,
         rowD_527,
         rowD_528,
         rowD_529,
         rowD_530,
         rowD_531,
         rowD_532,
         rowD_533,
         rowD_534,
         rowD_535,
         rowD_536,
         rowD_537,
         rowD_538,
         rowD_539,
         rowD_540,
         rowD_541,
         rowD_542,
         rowD_543,
         rowD_544,
         rowD_545,
         rowD_546,
         rowD_547,
         rowD_548,
         rowD_549,
         rowD_550,
         rowD_551,
         rowD_552,
         rowD_553,
         rowD_554,
         rowD_555,
         rowD_556,
         rowD_557,
         rowD_558,
         rowD_559,
         rowD_560,
         rowD_561,
         rowD_562,
         rowD_563,
         rowD_564,
         rowD_565,
         rowD_566,
         rowD_567,
         rowD_568,
         rowD_569,
         rowD_570,
         rowD_571,
         rowD_572,
         rowD_573,
         rowD_574,
         rowD_575,
         rowD_576,
         rowD_577,
         rowD_578,
         rowD_579,
         rowD_580,
         rowD_581,
         rowD_582,
         rowD_583,
         rowD_584,
         rowD_585,
         rowD_586,
         rowD_587,
         rowD_588,
         rowD_589,
         rowD_590,
         rowD_591,
         rowD_592,
         rowD_593,
         rowD_594,
         rowD_595,
         rowD_596,
         rowD_597,
         rowD_598,
         rowD_599,
         rowD_600,
         rowD_601,
         rowD_602,
         rowD_603,
         rowD_604,
         rowD_605,
         rowD_606,
         rowD_607,
         rowD_608,
         rowD_609,
         rowD_610,
         rowD_611,
         rowD_612,
         rowD_613,
         rowD_614,
         rowD_615,
         rowD_616,
         rowD_617,
         rowD_618,
         rowD_619,
         rowD_620,
         rowD_621,
         rowD_622,
         rowD_623,
         rowD_624,
         rowD_625,
         rowD_626,
         rowD_627,
         rowD_628,
         rowD_629,
         rowD_630,
         rowD_631,
         rowD_632,
         rowD_633,
         rowD_634,
         rowD_635,
         rowD_636,
         rowD_637,
         rowD_638,
         rowD_639,
         enP2S,
         ce_out4,
         pixel_out,
         enout
);  

endmodule
